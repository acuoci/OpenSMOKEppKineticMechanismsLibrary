! 
! CRECK Modeling Group (Politecnico di Milano)
! http://creckmodeling.chem.polimi.it/
! Version 1311, November 2013
!
 THERMO
  300.   1000.   4000.
HE                      HE  1               G    300.00   4000.00 1000.00      1
 .250000000E+01 .000000000E+00 .000000000E+00 .000000000E+00 .000000000E+00    2
-.745375000E+03 .928723974E+00 .250000000E+01 .000000000E+00 .000000000E+00    3
 .000000000E+00 .000000000E+00-.745375000E+03 .928723974E+00                   4
AR                      AR  1               G    300.00   4000.00 1000.00      1
 .250000000E+01 .000000000E+00 .000000000E+00 .000000000E+00 .000000000E+00    2
-.745375000E+03 .436600000E+01 .250000000E+01 .000000000E+00 .000000000E+00    3
 .000000000E+00 .000000000E+00-.745375000E+03 .436600000E+01                   4
N2                      N   2               G    300.00   4000.00 1000.00      1
 .292663788E+01 .148797700E-02-.568476030E-06 .100970400E-09-.675335090E-14    2
-.922795384E+03 .598054018E+01 .329867700E+01 .140823990E-02-.396322180E-05    3
 .564151480E-08-.244485400E-11-.102090000E+04 .395037200E+01                   4
NO                      O   1N   1          G    300.00   4000.00 1000.00      1
 .324543589E+01 .126913800E-02-.501589000E-06 .916928270E-10-.627541890E-14    2
 .980084032E+04 .641728767E+01 .337654100E+01 .125306300E-02-.330275000E-05    3
 .521781020E-08-.244626190E-11 .981796100E+04 .582959200E+01                   4
N2O                     O   1N   2          G    300.00   4000.00 1000.00      1
 .471897567E+01 .287371290E-02-.119749600E-05 .225055100E-09-.157533690E-13    2
 .816581343E+04-.165723704E+01 .254305700E+01 .949219330E-02-.979277500E-05    3
 .626384410E-08-.190182510E-11 .876510200E+04 .951122400E+01                   4
O2                      O   2               G    300.00   4000.00 1000.00      1
 .369757685E+01 .613519690E-03-.125884200E-06 .177528100E-10-.113643500E-14    2
-.123392966E+04 .318917125E+01 .321293600E+01 .112748610E-02-.575614990E-06    3
 .131387700E-08-.876855390E-12-.100524900E+04 .603473900E+01                   4
NO2                     O   2N   1          G    300.00   4000.00 1000.00      1
 .468285677E+01 .246242900E-02-.104225900E-05 .197690200E-09-.139171700E-13    2
 .226129300E+04 .988610659E+00 .267060000E+01 .783849970E-02-.806386380E-05    3
 .616171380E-08-.232014990E-11 .289629000E+04 .116120700E+02                   4
HNO                     H   1O   1N   1     G    300.00   4000.00 1000.00      1
 .361514436E+01 .321248500E-02-.126033690E-05 .226729700E-09-.153623600E-13    2
 .106619122E+05 .481025325E+01 .278440200E+01 .660964610E-02-.930022270E-05    3
 .943798020E-08-.375314580E-11 .109187800E+05 .903562900E+01                   4
HNNO                    H   1O   1N   2     G    300.00   4000.00 1500.00      1
 .699121930E+01 .187597000E-02-.212458400E-06-.671047200E-10 .123050800E-13    2
 .249756641E+05-.112352384E+02 .223829800E+01 .135920000E-01-.117987300E-04    3
 .539297100E-08-.101085900E-11 .266025900E+05 .141367900E+02                   4
HONO                    H   1O   2N   1     G    300.00   4000.00 1000.00      1
 .548688978E+01 .421806500E-02-.164914300E-05 .297187700E-09-.202114800E-13    2
-.112686489E+05-.299698546E+01 .229041300E+01 .140992200E-01-.136787200E-04    3
 .749878000E-08-.187690500E-11-.104319500E+05 .132807700E+02                   4
HNO2                    H   1O   2N   1     G    300.00   4000.00 1500.00      1
 .647962840E+01 .199527400E-02-.174038700E-06-.969587200E-10 .170148000E-13    2
-.999926943E+04-.106728455E+02 .193483800E+01 .101003600E-01-.496461600E-05    3
 .870112000E-09-.232413500E-14-.810548400E+04 .147325000E+02                   4
HONO2                   H   1O   3N   1     G    300.00   4000.00 1500.00      1
 .975613289E+01 .190094800E-02-.324002000E-06-.397663900E-10 .110033400E-13    2
-.194224157E+05-.269001236E+02 .787766800E+00 .238232900E-01-.220596400E-04    3
 .103404800E-07-.197285700E-11-.163044200E+05 .210896400E+02                   4
H2                      H   2               G    300.00   4000.00 1000.00      1
 .299142220E+01 .700064410E-03-.563382800E-07-.923157820E-11 .158275200E-14    2
-.835033546E+03-.135510641E+01 .329812400E+01 .824944120E-03-.814301470E-06    3
-.947543430E-10 .413487200E-12-.101252100E+04-.329409400E+01                   4
N2H2                    H   2N   2          G    300.00   4000.00 1000.00      1
 .337118994E+01 .603996800E-02-.230385300E-05 .406278900E-09-.271314400E-13    2
 .241817095E+05 .498055769E+01 .161799940E+01 .130631220E-01-.171571100E-04    3
 .160560790E-07-.609363800E-11 .246752600E+05 .137946700E+02                   4
H2O                     H   2O   1          G    300.00   4000.00 1000.00      1
 .267214569E+01 .305629290E-02-.873026070E-06 .120099600E-09-.639161790E-14    2
-.298992115E+05 .686281125E+01 .338684200E+01 .347498200E-02-.635469590E-05    3
 .696858040E-08-.250658800E-11-.302081100E+05 .259023200E+01                   4
H2O2                    H   2O   2          G    300.00   4000.00 1000.00      1
 .457316594E+01 .433613590E-02-.147468900E-05 .234890300E-09-.143165410E-13    2
-.180069531E+05 .501137915E+00 .338875300E+01 .656922580E-02-.148501200E-06    3
-.462580510E-08 .247151410E-11-.176631400E+05 .678536300E+01                   4
NH3                     H   3N   1          G    300.00   4000.00 1000.00      1
 .246189456E+01 .605916650E-02-.200497610E-05 .313600310E-09-.193831700E-13    2
-.649326483E+04 .747215046E+01 .220435100E+01 .101147600E-01-.146526500E-04    3
 .144723500E-07-.532850890E-11-.652548900E+04 .812714000E+01                   4
N2H4                    H   4N   2          G    300.00   4000.00 1000.00      1
 .497732211E+01 .959551900E-02-.354763900E-05 .612429900E-09-.402979500E-13    2
 .934121983E+04-.296302077E+01 .644260600E-01 .274973000E-01-.289945100E-04    3
 .174524000E-07-.442228200E-11 .104519200E+05 .212778900E+02                   4
CO                      C   1O   1          G    300.00   4000.00 1000.00      1
 .302507617E+01 .144268900E-02-.563082720E-06 .101858100E-09-.691095110E-14    2
-.142683499E+05 .610822521E+01 .326245100E+01 .151194100E-02-.388175520E-05    3
 .558194380E-08-.247495100E-11-.143105400E+05 .484889700E+01                   4
CO2                     C   1O   2          G    300.00   4000.00 1000.00      1
 .445362582E+01 .314016800E-02-.127841100E-05 .239399610E-09-.166903300E-13    2
-.489669524E+05-.955420007E+00 .227572400E+01 .992207230E-02-.104091100E-04    3
 .686668590E-08-.211728010E-11-.483731400E+05 .101884900E+02                   4
HCN                     C   1H   1N   1     G    300.00   4000.00 1000.00      1
 .365007798E+01 .346099790E-02-.127427900E-05 .221765490E-09-.147717700E-13    2
 .149839102E+05 .239321426E+01 .249046200E+01 .861127950E-02-.103103400E-04    3
 .748149810E-08-.222910900E-11 .152083400E+05 .790498000E+01                   4
HOCN                    C   1H   1O   1N   1G    300.00   4000.00 1000.00      1
 .564560836E+01 .229820610E-02-.216262900E-06-.121480100E-09 .223863610E-13    2
-.317811025E+04-.359027798E+01 .362829200E+01 .566418420E-02-.117020600E-06    3
-.234863800E-08 .801640220E-12-.247592500E+04 .747682300E+01                   4
HCNO                    C   1H   1O   1N   1G    300.00   4000.00 1000.00      1
 .669241213E+01 .236836030E-02-.237151000E-06-.127550300E-09 .240713700E-13    2
 .169473623E+05-.124543537E+02 .318485800E+01 .975231640E-02-.128020300E-05    3
-.616310380E-08 .322627490E-11 .179790700E+05 .612384200E+01                   4
HNCO                    C   1H   1O   1N   1G    300.00   4000.00 1000.00      1
 .621186395E+01 .229713690E-02-.221612790E-06-.122204400E-09 .227240590E-13    2
-.147707257E+05-.801661658E+01 .369405900E+01 .665723530E-02-.505446810E-07    3
-.347341090E-08 .136056900E-11-.139197600E+05 .571273900E+01                   4
CH2O                    C   1H   2O   1     G    300.00   4000.00 1000.00      1
 .299560858E+01 .668132120E-02-.262895400E-05 .473715290E-09-.321251710E-13    2
-.153203666E+05 .691256052E+01 .165273100E+01 .126314400E-01-.188816790E-04    3
 .205003110E-07-.841323710E-11-.148654000E+05 .137848200E+02                   4
HCOOH                   C   1H   2O   2     G    300.00   4000.00 1376.00      1
 .668733013E+01 .514289368E-02-.182238513E-05 .289719163E-09-.170892199E-13    2
-.483995400E+05-.113104798E+02 .143548185E+01 .163363016E-01-.106257421E-04    3
 .332132977E-08-.402176103E-12-.464616504E+05 .172885798E+02                   4
HCO3H                   C   1H   2O   3     G    300.00   4000.00 1378.00      1
 .987503581E+01 .464663708E-02-.167230522E-05 .268624413E-09-.159595232E-13    2
-.380502456E+05-.224938942E+02 .242464726E+01 .219706380E-01-.168705546E-04    3
 .625612194E-08-.911645843E-12-.354828006E+05 .175027796E+02                   4
CH3NO                   C   1H   3O   1N   1G    300.00   4000.00 1500.00      1
 .882055478E+01 .370623300E-02-.289474100E-06-.189791000E-09 .323754400E-13    2
 .536285603E+04-.221322539E+02 .210995500E+01 .151782200E-01-.707178900E-05    3
 .151061100E-08-.160420400E-12 .829361200E+04 .156970200E+02                   4
CH3ONO                  C   1H   3O   2N   1G    300.00   4000.00 1500.00      1
 .113612738E+02 .415934900E-02-.414567000E-06-.169514000E-09 .302873200E-13    2
-.128147952E+05-.354542296E+02 .149034500E+01 .264543300E-01-.211233200E-04    3
 .941439900E-08-.181120500E-11-.912578200E+04 .181376600E+02                   4
CH3NO2                  C   1H   3O   2N   1G    300.00   4000.00 1382.00      1
 .750407068E+01 .952121946E-02-.327760562E-05 .508678596E-09-.294455378E-13    2
-.121591399E+05-.115088778E+02-.370775080E+00 .283702793E-01-.208339624E-04    3
 .808980673E-08-.130521082E-11-.945681543E+04 .306459151E+02                   4
CH3ONO2                 C   1H   3O   3N   1G    300.00   4000.00 1500.00      1
 .143618741E+02 .411224300E-02-.511305200E-06-.149643600E-09 .301215600E-13    2
-.197243835E+05-.513183467E+02 .780335400E+00 .345420400E-01-.282232800E-04    3
 .123232400E-07-.230216400E-11-.146534600E+05 .224575200E+02                   4
CH4                     C   1H   4          G    300.00   4000.00 1000.00      1
 .168346564E+01 .102372400E-01-.387512820E-05 .678558490E-09-.450342310E-13    2
-.100807773E+05 .962347575E+01 .778741700E+00 .174766800E-01-.278340900E-04    3
 .304970800E-07-.122393100E-10-.982522800E+04 .137221900E+02                   4
CH3OH                   C   1H   4O   1     G    300.00   4000.00 1000.00      1
 .402907793E+01 .937659290E-02-.305025380E-05 .435879300E-09-.222472310E-13    2
-.261579223E+05 .237808255E+01 .266011500E+01 .734150780E-02 .717005010E-05    3
-.879319370E-08 .239056990E-11-.253534800E+05 .112326300E+02                   4
CH3OOH                  C   1H   4O   2     G    300.00   4000.00 1000.00      1
 .563694993E+01 .111814780E-01-.369593390E-05 .407189810E-09 .000000000E+00    2
-.180442749E+05-.124166637E+01 .586865100E+01 .107942400E-01-.364552990E-05    3
 .541291180E-09-.289684390E-13-.181268900E+05-.251762300E+01                   4
C2H2                    C   2H   2          G    300.00   4000.00 1000.00      1
 .443677300E+01 .537603910E-02-.191281610E-05 .328637890E-09-.215670900E-13    2
 .256676622E+05-.280035722E+01 .201356200E+01 .151904500E-01-.161631910E-04    3
 .907899180E-08-.191274600E-11 .261244400E+05 .880537800E+01                   4
CH2CO                   C   2H   2O   1     G    300.00   4000.00 1000.00      1
 .603885318E+01 .580484000E-02-.192095400E-05 .279448500E-09-.145886800E-13    2
-.858343402E+04-.765782305E+01 .297497100E+01 .121187100E-01-.234504600E-05    3
-.646668500E-08 .390564900E-11-.763263700E+04 .867355300E+01                   4
C2H2O2                  C   2H   2O   2     G    300.00   4000.00 1386.00      1
 .975438561E+01 .497645947E-02-.174410483E-05 .275586994E-09-.161969892E-13    2
-.295832896E+05-.261878329E+02 .188105120E+01 .236386368E-01-.183443295E-04    3
 .684842963E-08-.992733674E-12-.269280190E+05 .159154793E+02                   4
CH3CN                   C   2H   3N   1     G    300.00   4000.00 1000.00      1
 .239240386E+01 .156188730E-01-.791204970E-05 .193723330E-08-.186119560E-12    2
 .849993803E+04 .111452402E+02 .251975310E+01 .135675230E-01-.257640770E-05    3
-.308939670E-08 .142886920E-11 .855337620E+04 .109208680E+02                   4
C2H4                    C   2H   4          G    300.00   4000.00 1000.00      1
 .352841648E+01 .114851800E-01-.441838480E-05 .784460000E-09-.526684780E-13    2
 .442829030E+04 .223039249E+01-.861487900E+00 .279616190E-01-.338867690E-04    3
 .278515200E-07-.973787890E-11 .557304700E+04 .242114800E+02                   4
CH3CHO                  C   2H   4O   1     G    300.00   4000.00 1000.00      1
 .586869116E+01 .107942400E-01-.364552990E-05 .541291180E-09-.289684390E-13    2
-.226457128E+05-.601321650E+01 .250569500E+01 .133699100E-01 .467195290E-05    3
-.112814000E-07 .426356610E-11-.212458800E+05 .133508900E+02                   4
C2H4O                   C   2H   4O   1     G    300.00   4000.00 1000.00      1
 .385543260E+01 .146081760E-01-.526121540E-05 .628115500E-09 .000000000E+00    2
-.851874300E+04 .214156911E+01-.130385500E+01 .282461720E-01-.170593430E-04    3
 .394753470E-08 .000000000E+00-.707559900E+04 .289352600E+02                   4
CH3OCHO                 C   2H   4O   2     G    300.00   4000.00 1686.00      1
 .869123518E+01 .115503122E-01-.427782486E-05 .702533059E-09-.424333552E-13    2
-.464364769E+05-.189301478E+02 .308839783E+01 .203760048E-01-.684777040E-05    3
-.728186203E-09 .562130216E-12-.441855167E+05 .125364719E+02                   4
C2H4O2                  C   2H   4O   2     G    300.00   4000.00 1358.00      1
 .887306567E+01 .992257253E-02-.334820779E-05 .515546009E-09-.297527820E-13    2
-.410084739E+05-.182786314E+02 .437688685E+01 .159485358E-01-.363672718E-05    3
-.179212805E-08 .741898956E-12-.389689472E+05 .750888268E+01                   4
CH3COOH                 C   2H   4O   2     G    300.00   4000.00 1000.00      1
 .691666936E+01 .128920800E-01-.420990320E-05 .458049540E-09 .000000000E+00    2
-.553508487E+05-.102392103E+02 .846928500E+00 .292145000E-01-.186455200E-04    3
 .464098720E-08 .000000000E+00-.536761800E+05 .211901500E+02                   4
C2-OQOOH                C   2H   4O   3     G    300.00   4000.00 1380.00      1
 .124064339E+02 .947233784E-02-.328107928E-05 .513772211E-09-.299872803E-13    2
-.349123142E+05-.339479874E+02 .552382546E+01 .242068306E-01-.152898974E-04    3
 .501728362E-08-.696406358E-12-.323406789E+05 .357240645E+01                   4
CH3CO3H                 C   2H   4O   3     G    300.00   4000.00 1000.00      1
 .114777196E+02 .831667150E-02-.185084560E-05 .103274160E-09 .000000000E+00    2
-.451075908E+05-.290204723E+02 .484746000E+01 .218580610E-01-.904284660E-05    3
 .384145300E-09 .000000000E+00-.429209100E+05 .674072600E+01                   4
DME-OQOOH               C   2H   4O   4     G    300.00   4000.00 1000.00      1
 .114777196E+02 .831667150E-02-.185084560E-05 .103274160E-09 .000000000E+00    2
-.451075908E+05-.290204723E+02 .484746000E+01 .218580610E-01-.904284660E-05    3
 .384145300E-09 .000000000E+00-.429209100E+05 .674072600E+01                   4
C2H6                    C   2H   6          G    300.00   4000.00 1000.00      1
 .482597579E+01 .138404300E-01-.455725790E-05 .672496720E-09-.359816110E-13    2
-.127178296E+05-.523976258E+01 .146253900E+01 .154946700E-01 .578050690E-05    3
-.125783200E-07 .458626710E-11-.112391800E+05 .144322900E+02                   4
CH3OCH3                 C   2H   6O   1     G    300.00   4000.00 1368.00      1
 .827732656E+01 .132135539E-01-.453264362E-05 .705316507E-09-.409933283E-13    2
-.261980897E+05-.215181376E+02 .150763450E+01 .239914228E-01-.868910500E-05    3
-.966835762E-10 .489319361E-12-.232810894E+05 .167317297E+02                   4
C2H5OH                  C   2H   6O   1     G    300.00   4000.00 1000.00      1
 .434717120E+01 .186288000E-01-.677946700E-05 .816592600E-09 .000000000E+00    2
-.306615743E+05 .324247304E+01 .576535800E+00 .289451200E-01-.161002000E-04    3
 .359164100E-08 .000000000E+00-.296359500E+05 .227081300E+02                   4
C2H5OOH                 C   2H   6O   2     G    300.00   4000.00 1000.00      1
 .914611907E+01 .144611400E-01-.455120020E-05 .475780030E-09 .000000000E+00    2
-.236690607E+05-.205899250E+02 .223998300E+01 .310914290E-01-.170933710E-04    3
 .329379790E-08 .000000000E+00-.216018500E+05 .158174300E+02                   4
GLIET                   C   2H   6O   2     G    300.00   4000.00 1401.00      1
 .936137341E+01 .139727496E-01-.460325193E-05 .696470779E-09-.396758376E-13    2
-.507704265E+05-.211659058E+02 .875442184E+00 .347430045E-01-.244109224E-04    3
 .942412745E-08-.152824605E-11-.479084203E+05 .240879974E+02                   4
C3H2                    C   3H   2          G    300.00   4000.00 1000.00      1
 .767099642E+01 .274874900E-02-.437094300E-06-.645559900E-10 .166388700E-13    2
 .625972092E+05-.123689926E+02 .316671400E+01 .248257200E-01-.459163700E-04    3
 .426801900E-07-.148215200E-10 .635042100E+05 .886944600E+01                   4
PC3H4                   C   3H   4          G    300.00   4000.00 1000.00      1
 .281460543E+01 .185524496E-01-.955026768E-05 .239951370E-08-.237485257E-12    2
 .207010771E+05 .860604972E+01 .146175323E+01 .246026602E-01-.190219395E-04    3
 .860363422E-08-.166729240E-11 .209209793E+05 .149262585E+02                   4
AC3H4                   C   3H   4          G    300.00   4000.00 1400.07      1
 .977625145E+01 .530213820E-02-.370111790E-06-.302638610E-09 .508958110E-13    2
 .195497314E+05-.307705909E+02 .253983090E+01 .163343700E-01-.176495000E-05    3
-.464736520E-08 .172913110E-11 .225124300E+05 .993570230E+01                   4
C2H3CHO                 C   3H   4O   1     G    300.00   4000.00 1393.00      1
 .104184607E+02 .948963321E-02-.329310529E-05 .516279203E-09-.301587291E-13    2
-.149629790E+05-.307232511E+02 .292355162E+00 .354321417E-01-.294936324E-04    3
 .128100124E-07-.226144108E-11-.116521584E+05 .228878280E+02                   4
C3H4O2                  C   3H   4O   2     G    300.00   4000.00 1404.00      1
 .130577477E+02 .906905120E-02-.308189261E-05 .476481380E-09-.275669277E-13    2
-.369274825E+05-.425273740E+02 .147485987E+00 .464706296E-01-.451901760E-04    3
 .219641008E-07-.416219125E-11-.331809255E+05 .242182934E+02                   4
C3H4O3                  C   3H   4O   3     G    300.00   4000.00 1388.00      1
 .137530675E+02 .108054207E-01-.364230159E-05 .560730953E-09-.323659923E-13    2
-.577839662E+05-.401019465E+02 .208981535E+01 .383715226E-01-.282590499E-04    3
 .104299134E-07-.153140407E-11-.538199819E+05 .223338530E+02                   4
C3H6                    C   3H   6          G    300.00   4000.00 1000.00      1
 .673231663E+01 .149083400E-01-.494989900E-05 .721202210E-09-.376620390E-13    2
-.923623057E+03-.133137684E+02 .149330700E+01 .209251700E-01 .448679380E-05    3
-.166891190E-07 .715814600E-11 .107482600E+04 .161453400E+02                   4
C3H6O                   C   3H   6O   1     G    300.00   4000.00 1000.00      1
 .433142310E+01 .236433890E-01-.875060690E-05 .106889830E-08 .000000000E+00    2
-.138496111E+05 .215169726E+01 .507423500E+00 .318789710E-01-.137497700E-04    3
 .165647900E-08 .000000000E+00-.126239100E+05 .226350900E+02                   4
CH3COCH3                C   3H   6O   1     G    300.00   4000.00 1374.00      1
 .991426580E+01 .146030709E-01-.506085765E-05 .792682855E-09-.462739645E-13    2
-.311168055E+05-.286116537E+02 .130767163E+01 .292021742E-01-.119045617E-04    3
 .652150087E-09 .467751203E-12-.275328269E+05 .196395025E+02                   4
C3H5OH                  C   3H   6O   1     G    300.00   4000.00 1000.00      1
 .665875100E+01 .179008100E-01-.612801520E-05 .983706560E-09-.609475850E-13    2
-.187194550E+05-.446185680E+01 .332545570E+01 .251539630E-01-.163055650E-04    3
 .121609030E-07-.500807290E-11-.174250940E+05 .139104030E+02                   4
C2H5CHO                 C   3H   6O   1     G    300.00   4000.00 1378.00      1
 .102429148E+02 .139641989E-01-.476248001E-05 .738105706E-09-.427759503E-13    2
-.274145137E+05-.285357348E+02 .216308444E+01 .295501264E-01-.152446252E-04    3
 .349503947E-08-.238896627E-12-.242260137E+05 .161153348E+02                   4
C3H5OOH                 C   3H   6O   2     G    300.00   4000.00 1382.00      1
 .139268456E+02 .135384067E-01-.474335693E-05 .748389157E-09-.439105886E-13    2
-.132537727E+05-.456757848E+02 .221491505E+01 .390935107E-01-.258809564E-04    3
 .870894601E-08-.120793929E-11-.896037969E+04 .179425329E+02                   4
C3H6O2                  C   3H   6O   2     G    300.00   4000.00 1382.00      1
 .118936666E+02 .144153203E-01-.477525443E-05 .726036430E-09-.415285995E-13    2
-.459271652E+05-.327285750E+02 .266613285E+01 .346302298E-01-.214380719E-04    3
 .690469334E-08-.916939105E-12-.425706030E+05 .173358364E+02                   4
ACETOL                  C   3H   6O   2     G    300.00   4000.00 1390.00      1
 .110277409E+02 .156022896E-01-.518498789E-05 .789604263E-09-.452017356E-13    2
-.493518932E+05-.296460029E+02 .170110573E+01 .349995386E-01-.195672111E-04    3
 .513929120E-08-.454830190E-12-.458857790E+05 .212715964E+02                   4
C3-OQOOH                C   3H   6O   3     G    300.00   4000.00 1391.00      1
 .170285271E+02 .130716784E-01-.459310856E-05 .726135156E-09-.426658337E-13    2
-.416334217E+05-.592513577E+02 .768933034E+00 .546905880E-01-.465072405E-04    3
 .203159585E-07-.358398999E-11-.363238861E+05 .268291637E+02                   4
C3H8                    C   3H   8          G    300.00   4000.00 1000.00      1
 .752530602E+01 .188903400E-01-.628392400E-05 .917937280E-09-.481240960E-13    2
-.164646226E+05-.178445202E+02 .896921000E+00 .266898590E-01 .543142510E-05    3
-.212600000E-07 .924333010E-11-.139549200E+05 .193553300E+02                   4
IC3H7OH                 C   3H   8O   1     G    300.00   4000.00 1000.00      1
 .577239007E+01 .268947430E-01-.111795290E-04 .211392460E-08-.149320990E-12    2
-.361710675E+05-.384089810E+01-.176838920E+00 .452559560E-01-.319190720E-04    3
 .123062880E-07-.201412540E-11-.346643940E+05 .263322250E+02                   4
NC3H7OH                 C   3H   8O   1     G    300.00   4000.00 1396.00      1
 .107520626E+02 .180260472E-01-.603049401E-05 .922166246E-09-.529319319E-13    2
-.361555719E+05-.310977038E+02 .978207214E-01 .420500918E-01-.267066894E-04    3
 .903941170E-08-.128324751E-11-.323437836E+05 .264700804E+02                   4
C3H7OOH                 C   3H   8O   2     G    300.00   4000.00 1388.00      1
 .150655849E+02 .170865595E-01-.593183927E-05 .930136673E-09-.543384935E-13    2
-.301371140E+05-.515057998E+02 .783525746E+00 .504826223E-01-.365089942E-04    3
 .140377750E-07-.226737156E-11-.251105573E+05 .253041175E+02                   4
GLYCEROL                C   3H   8O   3     G    300.00   4000.00 1413.00      1
 .142234482E+02 .188282751E-01-.593875071E-05 .871197709E-09-.485331087E-13    2
-.753882525E+05-.411276527E+02 .214180274E+00 .584817984E-01-.493063032E-04    3
 .223333179E-07-.405800253E-11-.712682818E+05 .315639747E+02                   4
C4H2                    C   4H   2          G    300.00   4000.00 1000.00      1
 .903147468E+01 .604725210E-02-.194878790E-05 .275486300E-09-.138560800E-13    2
 .529472934E+05-.238511290E+02 .400519100E+01 .198100000E-01-.986587660E-05    3
-.663515820E-08 .607741290E-11 .542406400E+05 .184573600E+01                   4
C4H4                    C   4H   4          G    300.00   4000.00 1000.00      1
 .665080310E+01 .161294300E-01-.719388700E-05 .149817800E-08-.118641100E-12    2
 .311958636E+05-.979559836E+01-.191524700E+01 .527508700E-01-.716559400E-04    3
 .550724200E-07-.172862200E-10 .329785000E+05 .314199800E+02                   4
C4H4O                   C   4H   4O   1     G    300.00   4000.00 1000.00      1
 .135912211E+02 .987450910E-02-.345325238E-05 .544429808E-09-.319349896E-13    2
-.115639534E+05-.542513644E+02-.750030326E+01 .699899868E-01-.695485649E-04    3
 .333968809E-07-.619467883E-11-.541634292E+04 .550218432E+02                   4
CH2CCHCHO               C   4H   4O   1     G    300.00   4000.00 1000.00      1
 .929991052E+01 .152201510E-01-.615883937E-05 .112678366E-08-.769359137E-13    2
 .368009609E+04-.220663746E+02 .123852148E+01 .356054647E-01-.236786887E-04    3
 .592234361E-08 .282885884E-12 .610569242E+04 .202911558E+02                   4
C4H6                    C   4H   6          G    300.00   4000.00 1000.00      1
 .823794980E+01 .173695890E-01-.615923200E-05 .979908060E-09-.578075590E-13    2
 .923259930E+04-.203418190E+02 .112443850E+00 .343711770E-01-.111106630E-04    3
-.921096660E-08 .620841700E-11 .118022620E+05 .230917180E+02                   4
IC3H5CHO                C   4H   6O   1     G    300.00   4000.00 1396.00      1
 .136175682E+02 .137917192E-01-.473370118E-05 .736655226E-09-.420097974E-13    2
-.199994281E+05-.472987367E+02 .627183793E+00 .466780254E-01-.374430631E-04    3
 .158330542E-07-.273952155E-11-.157203117E+05 .216034294E+02                   4
C4H6O2                  C   4H   6O   2     G    300.00   4000.00 1375.00      1
 .135393551E+02 .168328392E-01-.587873230E-05 .925553795E-09-.542254877E-13    2
-.462482008E+05-.437360830E+02 .182538964E+01 .377978336E-01-.172044878E-04    3
 .195698878E-08 .398612932E-12-.415126261E+05 .214925508E+02                   4
MACRIL                  C   4H   6O   2     G    300.00   4000.00 1000.00      1
 .962595080E+01 .202069860E-01-.684948550E-05 .109063620E-08-.671284990E-13    2
-.414857110E+05-.177414250E+02-.929250120E+00 .565245670E-01-.531143270E-04    3
 .263405850E-07-.484636380E-11-.390243280E+05 .347643170E+02                   4
NC4H8                   C   4H   8          G    300.00   4000.00 1000.00      1
 .205358410E+01 .343505070E-01-.158831970E-04 .330896620E-08-.253610450E-12    2
-.213972310E+04 .155432010E+02 .118113800E+01 .308533800E-01 .508652470E-05    3
-.246548880E-07 .111101930E-10-.179040040E+04 .210624690E+02                   4
IC4H8                   C   4H   8          G    300.00   4000.00 1388.00      1
 .112258330E+02 .181795798E-01-.620348592E-05 .961444458E-09-.557088057E-13    2
-.769983777E+04-.373306704E+02 .938433173E+00 .390547287E-01-.216437148E-04    3
 .587267077E-08-.614435479E-12-.374817891E+04 .191442985E+02                   4
C4H8O                   C   4H   8O   1     G    300.00   4000.00 1371.00      1
 .154228514E+02 .170211052E-01-.606347951E-05 .967354762E-09-.571992419E-13    2
-.220196123E+05-.613882135E+02-.253690104E+01 .543995707E-01-.343390305E-04    3
 .101079922E-07-.110262736E-11-.152980680E+05 .367400719E+02                   4
MEK                     C   4H   8O   1     G    300.00   4000.00 1000.00      1
 .929655016E+01 .229172746E-01-.822048591E-05 .132404838E-08-.791751980E-13    2
-.334442311E+05-.204993263E+02 .661978185E+01 .851847835E-02 .510322077E-04    3
-.658433042E-07 .249110484E-10-.315251691E+05-.109485469E+01                   4
C4H7OH                  C   4H   8O   1     G    300.00   4000.00 1000.00      1
 .863167950E+01 .241150480E-01-.832957180E-05 .134433130E-08-.835340300E-13    2
-.230779140E+05-.163015210E+02 .173864090E+01 .369849060E-01-.680297030E-05    3
-.128647340E-07 .662652570E-11-.209184180E+05 .207395880E+02                   4
C3H7CHO                 C   4H   8O   1     G    300.00   4000.00 1000.00      1
 .885754490E+01 .242627260E-01-.846559850E-05 .137561310E-08-.858588980E-13    2
-.294816840E+05-.174775160E+02 .666312930E+00 .477311800E-01-.329931100E-04    3
 .121733550E-07-.165405020E-11-.272346390E+05 .246936170E+02                   4
IC3H7CHO                C   4H   8O   1     G    300.00   4000.00 1391.00      1
 .137503148E+02 .183126722E-01-.628572629E-05 .978250756E-09-.568538653E-13    2
-.326938845E+05-.477281342E+02-.273021382E+00 .489696307E-01-.312770049E-04    3
 .100052945E-07-.127512074E-11-.276054737E+05 .283451139E+02                   4
NC4-OQOOH               C   4H   8O   3     G    300.00   4000.00 1388.00      1
 .195955254E+02 .180568312E-01-.629994700E-05 .991157547E-09-.580382406E-13    2
-.461054913E+05-.709333761E+02 .243440296E+01 .605409309E-01-.481250984E-04    3
 .203656751E-07-.357059537E-11-.402872220E+05 .205488821E+02                   4
IC4-OQOOH               C   4H   8O   3     G    300.00   4000.00 1390.00      1
 .195047991E+02 .181701803E-01-.634838146E-05 .999797067E-09-.585883751E-13    2
-.450007951E+05-.705122130E+02 .549934041E+00 .642751153E-01-.501779820E-04    3
 .203546231E-07-.338767418E-11-.385647626E+05 .307013051E+02                   4
KEHYBU1                 C   4H   8O   4     G    300.00   4000.00 1396.00      1
 .219367270E+02 .180406285E-01-.626171080E-05 .981855896E-09-.573639516E-13    2
-.664546784E+05-.813588272E+02-.445736457E+01 .947202096E-01-.937478682E-04    3
 .464802131E-07-.899314409E-11-.587131282E+05 .551970961E+02                   4
NC4H10                  C   4H  10          G    300.00   4000.00 1000.00      1
 .105251152E+02 .235908740E-01-.785389060E-05 .114561140E-08-.599309560E-13    2
-.204952316E+05-.321928008E+02 .157641510E+01 .345897230E-01 .697016090E-05    3
-.281636370E-07 .123751170E-10-.171470040E+05 .178727420E+02                   4
IC4H10                  C   4H  10          G    300.00   4000.00 1000.00      1
 .508434390E+01 .331851280E-01-.124047670E-04 .152753620E-08 .000000000E+00    2
-.195243797E+05-.392308050E+01-.128398800E+01 .519486400E-01-.308267920E-04    3
 .755438110E-08 .000000000E+00-.179038400E+05 .285063500E+02                   4
N2C4H9OH                C   4H  10O   1     G    300.00   4000.00 1390.00      1
 .151582366E+02 .215048627E-01-.741631184E-05 .115764678E-08-.674130532E-13    2
-.429113728E+05-.549620416E+02-.304705097E+00 .567446943E-01-.387293873E-04    3
 .141775813E-07-.220696859E-11-.373601662E+05 .285520284E+02                   4
TC4H9OH                 C   4H  10O   1     G    300.00   4000.00 1395.00      1
 .151183592E+02 .214941230E-01-.730928419E-05 .113021881E-08-.653833962E-13    2
-.450124898E+05-.575375902E+02-.861795957E+00 .603867730E-01-.445191256E-04    3
 .177406426E-07-.295852901E-11-.395611057E+05 .278278048E+02                   4
N1C4H9OH                C   4H  10O   1     G    300.00   4000.00 1389.00      1
 .146461472E+02 .217370421E-01-.745243572E-05 .115877769E-08-.672987557E-13    2
-.406432319E+05-.509926617E+02 .129085275E+00 .529074664E-01-.325907761E-04    3
 .102723019E-07-.133027252E-11-.352672374E+05 .280463660E+02                   4
IC4H9OH                 C   4H  10O   1     G    300.00   4000.00 1426.00      1
 .145203606E+02 .218826590E-01-.741886985E-05 .114493281E-08-.661481541E-13    2
-.415815847E+05-.516504190E+02-.808654483E+00 .568695746E-01-.379891888E-04    3
 .133635469E-07-.195588405E-11-.361485459E+05 .310126347E+02                   4
C4H9OOH                 C   4H  10O   2     G    300.00   4000.00 1389.00      1
 .182257559E+02 .215996217E-01-.748424942E-05 .117205153E-08-.684096331E-13    2
-.342341151E+05-.670536388E+02 .607792497E+00 .624669916E-01-.444490375E-04    3
 .167754668E-07-.265938189E-11-.280070327E+05 .278025473E+02                   4
CYC5H4O                 C   5H   4O   1     G    300.00   4000.00 1000.00      1
 .558734350E+01 .254149730E-01-.929145880E-05 .112347330E-08 .000000000E+00    2
 .339172461E+04-.552979995E+01-.427809100E+01 .546170700E-01-.380993520E-04    3
 .105947040E-07 .000000000E+00 .589093400E+04 .446629800E+02                   4
C5H4O2                  C   5H   4O   2     G    300.00   4000.00 1000.00      1
 .159553578E+02 .122096134E-01-.419491662E-05 .654219009E-09-.381060338E-13    2
-.255664634E+05-.596830465E+02-.186260023E+01 .570946426E-01-.476338594E-04    3
 .197949337E-07-.326585828E-11-.197873020E+05 .347179869E+02                   4
CYC5H6                  C   5H   6          G    300.00   4000.00 1000.00      1
 .230537462E+00 .409571826E-01-.241588958E-04 .679763480E-08-.736374421E-12    2
 .143779465E+05 .202551234E+02-.513691194E+01 .606953453E-01-.460552837E-04    3
 .128457201E-07 .741214852E-12 .153675713E+05 .461567559E+02                   4
MEFU2                   C   5H   6O   1     G    300.00   4000.00 1000.00      1
 .459933100E+01 .340025700E-01-.175181400E-04 .423464670E-08-.375757330E-12    2
-.129526080E+05 .466753790E+00-.284971730E+01 .552316440E-01-.365110720E-04    3
 .832948240E-08 .742313490E-12-.110344430E+05 .385458850E+02                   4
CYC5H8                  C   5H   8          G    300.00   4000.00 1000.00      1
 .772447728E+01 .283223160E-01-.115452360E-04 .215408150E-08-.150541780E-12    2
-.782614232E+03-.197696844E+02 .268981400E+01 .209545500E-02 .113036870E-03    3
-.154080700E-06 .627636580E-10 .231396630E+04 .152940560E+02                   4
C5H8                    C   5H   8          G    300.00   4000.00 1000.00      1
 .797205310E+01 .268614160E-01-.956546320E-05 .113079120E-08 .000000000E+00    2
 .510466811E+04-.185090870E+02 .176636500E+01 .432678800E-01-.237613290E-04    3
 .512588110E-08 .000000000E+00 .684030700E+04 .137180600E+02                   4
C5H8O                   C   5H   8O   1     G    300.00   4000.00 1000.00      1
 .154011002E+02 .203490440E-01-.699742510E-05 .109031908E-08-.634192782E-13    2
-.910076428E+04-.580710041E+02-.514624016E+01 .722177875E-01-.580157542E-04    3
 .242093068E-07-.410120178E-11-.236133441E+04 .508920452E+02                   4
MCROT                   C   5H   8O   2     G    300.00   4000.00 1000.00      1
 .110840220E+02 .266681570E-01-.910298150E-05 .145819250E-08-.902072000E-13    2
-.461868520E+05-.238654710E+02 .115411390E+01 .550597160E-01-.356332020E-04    3
 .867407750E-08 .746845670E-12-.435806950E+05 .269868980E+02                   4
C5EN-OQOOH-53           C   5H   8O   3     G    300.00   4000.00 1389.00      1
 .217801959E+02 .189644170E-01-.666360530E-05 .105343196E-08-.618948648E-13    2
-.372541821E+05-.828559128E+02 .975948412E+00 .693438350E-01-.543693801E-04    3
 .220678107E-07-.367435527E-11-.301615960E+05 .283235620E+02                   4
ETMB583                 C   5H   8O   3     G    300.00   4000.00 1000.00      1
 .164044820E+02 .257082970E-01-.901921340E-05 .147114070E-08-.920586850E-13    2
-.622657890E+05-.550660710E+02-.249091940E+01 .790685040E-01-.564648800E-04    3
 .115540360E-07 .278656790E-11-.573317190E+05 .417407460E+02                   4
C5EN-OQOOH-54           C   5H   8O   3     G    300.00   4000.00 1389.00      1
 .217801959E+02 .189644170E-01-.666360530E-05 .105343196E-08-.618948648E-13    2
-.372541821E+05-.828559128E+02 .975948412E+00 .693438350E-01-.543693801E-04    3
 .220678107E-07-.367435527E-11-.301615960E+05 .283235620E+02                   4
C5EN-OQOOH-43           C   5H   8O   3     G    300.00   4000.00 1389.00      1
 .217801959E+02 .189644170E-01-.666360530E-05 .105343196E-08-.618948648E-13    2
-.372541821E+05-.828559128E+02 .975948412E+00 .693438350E-01-.543693801E-04    3
 .220678107E-07-.367435527E-11-.301615960E+05 .283235620E+02                   4
C5EN-OQOOH-45           C   5H   8O   3     G    300.00   4000.00 1389.00      1
 .217801959E+02 .189644170E-01-.666360530E-05 .105343196E-08-.618948648E-13    2
-.372541821E+05-.828559128E+02 .975948412E+00 .693438350E-01-.543693801E-04    3
 .220678107E-07-.367435527E-11-.301615960E+05 .283235620E+02                   4
C5EN-OQOOH-35           C   5H   8O   3     G    300.00   4000.00 1389.00      1
 .217801959E+02 .189644170E-01-.666360530E-05 .105343196E-08-.618948648E-13    2
-.372541821E+05-.828559128E+02 .975948412E+00 .693438350E-01-.543693801E-04    3
 .220678107E-07-.367435527E-11-.301615960E+05 .283235620E+02                   4
C5EN-OQOOH-34           C   5H   8O   3     G    300.00   4000.00 1389.00      1
 .217801959E+02 .189644170E-01-.666360530E-05 .105343196E-08-.618948648E-13    2
-.372541821E+05-.828559128E+02 .975948412E+00 .693438350E-01-.543693801E-04    3
 .220678107E-07-.367435527E-11-.301615960E+05 .283235620E+02                   4
C5H8O4                  C   5H   8O   4     G    300.00   4000.00 1000.00      1
 .217298154E+02 .217807665E-01-.749545594E-05 .116860895E-08-.680038942E-13    2
-.866505360E+05-.835752527E+02-.684199090E+01 .100610553E+00-.924172541E-04    3
 .429800586E-07-.789719358E-11-.779623201E+05 .655426910E+02                   4
KEHYMB                  C   5H   8O   5     G    300.00   4000.00 1000.00      1
 .130410150E+02 .302430520E-01-.103682550E-04 .166520830E-08-.103159200E-12    2
-.605793360E+05-.352927630E+02-.187604440E+01 .779613480E-01-.656695630E-04    3
 .280818550E-07-.405575270E-11-.569013010E+05 .398655930E+02                   4
IC5H10                  C   5H  10          G    300.00   4000.00 1000.00      1
 .124808598E+02 .240088830E-01-.777773490E-05 .119128510E-08-.709457860E-13    2
-.864177347E+04-.392940217E+02-.599261880E+00 .540460090E-01-.294562720E-04    3
 .525642110E-08 .585451010E-12-.450159910E+04 .303432560E+02                   4
NC5H10                  C   5H  10          G    300.00   4000.00 1389.00      1
 .141108203E+02 .228348272E-01-.778626835E-05 .120627491E-08-.698795983E-13    2
-.114335029E+05-.501593461E+02-.541560551E+00 .539629918E-01-.323508738E-04    3
 .977416037E-08-.118534668E-11-.598606169E+04 .297142748E+02                   4
NEOC5H10-O              C   5H  10O   1     G    300.00   4000.00 1406.00      1
 .182053093E+02 .222888126E-01-.759419141E-05 .117633164E-08-.681511068E-13    2
-.260973639E+05-.785614741E+02-.704702259E+01 .864172552E-01-.702610933E-04    3
 .290540959E-07-.480586102E-11-.179483330E+05 .550571499E+02                   4
NC5H10-O                C   5H  10O   1     G    300.00   4000.00 1373.00      1
 .187152768E+02 .216122625E-01-.768638433E-05 .122492227E-08-.723734176E-13    2
-.274341627E+05-.786690289E+02-.351633623E+01 .686975884E-01-.446579237E-04    3
 .140670556E-07-.174934766E-11-.191663581E+05 .425589840E+02                   4
C4H9CHO                 C   5H  10O   1     G    300.00   4000.00 1381.00      1
 .167965264E+02 .225684519E-01-.767631588E-05 .118769369E-08-.687545554E-13    2
-.356826220E+05-.609064044E+02 .159663472E+01 .543541416E-01-.321020651E-04    3
 .935773559E-08-.106688932E-11-.299841025E+05 .221281498E+02                   4
MB                      C   5H  10O   2     G    300.00   4000.00 1380.00      1
 .190094725E+02 .236503722E-01-.822978452E-05 .129246265E-08-.755862836E-13    2
-.634989152E+05-.732469099E+02 .316208825E+01 .552915358E-01-.311610102E-04    3
 .842394129E-08-.872222021E-12-.573385240E+05 .139723817E+02                   4
MTBE-O                  C   5H  10O   2     G    300.00   4000.00 1397.00      1
 .193844587E+02 .224929046E-01-.748169734E-05 .114123661E-08-.654437288E-13    2
-.558416627E+05-.795832532E+02-.518049059E+01 .839546669E-01-.663790553E-04    3
 .267623941E-07-.432034827E-11-.478415885E+05 .506953652E+02                   4
NC5-OQOOH               C   5H  10O   3     G    300.00   4000.00 1389.00      1
 .227422860E+02 .225948063E-01-.786379640E-05 .123514506E-08-.722413862E-13    2
-.501979972E+05-.864068664E+02 .227305950E+01 .724929431E-01-.560597536E-04    3
 .231254746E-07-.397203084E-11-.431866364E+05 .229745558E+02                   4
NEOC5-OQOOH             C   5H  10O   3     G    300.00   4000.00 1397.00      1
 .237028187E+02 .215843890E-01-.747470111E-05 .117038715E-08-.683143724E-13    2
-.509464263E+05-.948314143E+02 .101097520E+01 .753376897E-01-.559848192E-04    3
 .210040666E-07-.316727025E-11-.432003697E+05 .266737910E+02                   4
MTBE-OQOOH              C   5H  10O   4     G    300.00   4000.00 1386.00      1
 .259492704E+02 .217762181E-01-.754080079E-05 .118109778E-08-.689663912E-13    2
-.659884236E+05-.102260628E+03 .215705064E+01 .770950997E-01-.562944956E-04    3
 .205751475E-07-.301215733E-11-.577585957E+05 .255153989E+02                   4
NEOC5H12                C   5H  12          G    300.00   4000.00 1397.00      1
 .174488013E+02 .245462377E-01-.835182479E-05 .129219708E-08-.747942850E-13    2
-.292378530E+05-.754164601E+02-.288372771E+01 .722417687E-01-.511106166E-04    3
 .187342407E-07-.280628313E-11-.222171069E+05 .336765462E+02                   4
NC5H12                  C   5H  12          G    300.00   4000.00 1000.00      1
 .142233709E+02 .264253600E-01-.834599270E-05 .125651470E-08-.740004510E-13    2
-.247106388E+05-.503994927E+02-.393634560E+00 .578781330E-01-.285392090E-04    3
 .347472500E-08 .106523800E-11-.198713480E+05 .281908260E+02                   4
MTBE                    C   5H  12O   1     G    300.00   4000.00 1000.00      1
 .888656643E+01 .420057870E-01-.178904220E-04 .345077750E-08-.247674430E-12    2
-.405353691E+05-.208281992E+02-.162610860E+01 .742240170E-01-.539682020E-04    3
 .210023490E-07-.342702090E-11-.378579060E+05 .325557600E+02                   4
NC5H11OOH               C   5H  12O   2     G    300.00   4000.00 1391.00      1
 .215962451E+02 .259122865E-01-.896302814E-05 .140202940E-08-.817685827E-13    2
-.395542326E+05-.852046644E+02-.443227141E+00 .781363104E-01-.573273118E-04    3
 .222802059E-07-.361215684E-11-.318952281E+05 .330316890E+02                   4
C6H2                    C   6H   2          G    300.00   4000.00 1000.00      1
 .127565190E+02 .803438100E-02-.261821500E-05 .372506000E-09-.187885000E-13    2
 .807546900E+05-.404126200E+02 .575108500E+01 .263671900E-01-.116675960E-04    3
-.107144980E-07 .879029700E-11 .826201200E+05-.433553200E+01                   4
C6H4                    C   6H   4          G    300.00   4000.00 1000.00      1
 .171831170E+02 .664876580E-02-.124162630E-05 .146974480E-09-.913980130E-14    2
 .550769540E+05-.644351830E+02 .193231390E+01 .390321830E-01-.692271090E-05    3
-.270933570E-07 .157302520E-10 .596919480E+05 .165160230E+02                   4
BENZYNE                 C   6H   4          G    300.00   4000.00 1000.00      1
 .105707063E+02 .156860613E-01-.568267148E-05 .922956737E-09-.554966417E-13    2
 .504976657E+05-.332563927E+02 .721604591E+00 .247976151E-01 .316372209E-04    3
-.653230986E-07 .296082142E-10 .539797980E+05 .216733825E+02                   4
C6H4O2                  C   6H   4O   2     G    300.00   4000.00 1000.00      1
 .148186534E+02 .176963450E-01-.512229240E-05 .482867020E-09 .000000000E+00    2
-.210645982E+05-.499092297E+02-.357739600E+01 .669980650E-01-.485375860E-04    3
 .129924900E-07 .000000000E+00-.159750500E+05 .454022300E+02                   4
C6H6                    C   6H   6          G    300.00   4000.00 1000.00      1
 .129109067E+02 .172329600E-01-.502421020E-05 .589349680E-09-.194752100E-13    2
 .366437279E+04-.500281184E+02-.313801200E+01 .472310300E-01-.296220700E-05    3
-.326281900E-07 .171869100E-10 .889003000E+04 .365757300E+02                   4
LC6H6                   C   6H   6          G    300.00   4000.00 1000.00      1
 .133755312E+02 .181053970E-01-.671790940E-05 .114930710E-08-.753903640E-13    2
 .353349989E+05-.436278915E+02-.284372350E+01 .754240600E-01-.877316710E-04    3
 .551440390E-07-.141557690E-10 .392169020E+05 .371208190E+02                   4
C6H5OH                  C   6H   6O   1     G    300.00   4000.00 1000.00      1
 .141552427E+02 .199350340E-01-.718219540E-05 .116229002E-08-.697147483E-13    2
-.181287441E+05-.517984911E+02-.290978575E+00 .408562397E-01 .242829425E-04    3
-.714477617E-07 .346002146E-10-.134129780E+05 .268745637E+02                   4
C6H6O3                  C   6H   6O   3     G    300.00   4000.00 1382.00      1
 .193892545E+02 .186134462E-01-.631148097E-05 .975462374E-09-.564561412E-13    2
-.492678935E+05-.716786498E+02 .598814621E+00 .618493802E-01-.438009436E-04    3
 .155531333E-07-.220506530E-11-.427313109E+05 .293828012E+02                   4
CYC6H8                  C   6H   8          G    300.00   4000.00 1384.00      1
 .167797183E+02 .200748305E-01-.710732570E-05 .112925397E-08-.665827513E-13    2
 .222453062E+04-.729120687E+02-.719572313E+01 .780676798E-01-.620002183E-04    3
 .253310854E-07-.423684696E-11 .104082650E+05 .552451233E+02                   4
MCPTD                   C   6H   8          G    300.00   4000.00 1399.00      1
 .154352848E+02 .199801707E-01-.680270423E-05 .105349633E-08-.610336727E-13    2
 .447456576E+04-.636393642E+02-.665320026E+01 .744640477E-01-.582864186E-04    3
 .231603543E-07-.369017129E-11 .117669311E+05 .538162769E+02                   4
DMF                     C   6H   8O   1     G    300.00   4000.00 1000.00      1
 .117792073E+02 .285086757E-01-.111333319E-04 .199173491E-08-.133982691E-12    2
-.211130695E+05-.374257400E+02 .803526924E+00 .443305994E-01 .419434116E-05    3
-.349560898E-07 .165826978E-10-.172836857E+05 .230189579E+02                   4
C6H8O4                  C   6H   8O   4     G    300.00   4000.00 1398.00      1
 .245389912E+02 .222706283E-01-.773806446E-05 .121423501E-08-.709771757E-13    2
-.816610603E+05-.100550137E+03-.460104207E+01 .100736116E+00-.905484350E-04    3
 .413812870E-07-.752102026E-11-.725801173E+05 .522649333E+02                   4
CYC6H10                 C   6H  10          G    300.00   4000.00 1388.00      1
 .164687940E+02 .250464584E-01-.873323457E-05 .137353265E-08-.804138942E-13    2
-.977694533E+04-.696690108E+02-.607599781E+01 .751138370E-01-.506516889E-04    3
 .171683701E-07-.235089637E-11-.166592755E+04 .523699408E+02                   4
CYC6H10-O-12            C   6H  10O   1     G    300.00   4000.00 1388.00      1
 .211309516E+02 .245922161E-01-.870218393E-05 .138238722E-08-.815033630E-13    2
-.270082298E+05-.100017882E+03-.102441734E+02 .947119743E-01-.662992744E-04    3
 .218368996E-07-.269065692E-11-.159562249E+05 .693449458E+02                   4
C5H9CHO                 C   6H  10O   1     G    300.00   4000.00 1369.00      1
 .194648486E+02 .257619052E-01-.914519168E-05 .145563936E-08-.859339746E-13    2
-.393988116E+05-.858349504E+02-.528503736E+01 .742084262E-01-.414393902E-04    3
 .926068588E-08-.391839791E-12-.298547201E+05 .504370563E+02                   4
CYC6H10-O-14            C   6H  10O   1     G    300.00   4000.00 1381.00      1
 .208569012E+02 .251723586E-01-.898344923E-05 .143508332E-08-.849382249E-13    2
-.384586302E+05-.102070819E+03-.138345764E+02 .100994913E+00-.688346635E-04    3
 .212451763E-07-.229797219E-11-.260978348E+05 .857505804E+02                   4
CYC6H10-ONE             C   6H  10O   1     G    300.00   4000.00 1382.00      1
 .189587175E+02 .263606964E-01-.929344737E-05 .147257311E-08-.866645349E-13    2
-.391424596E+05-.835594309E+02-.541298687E+01 .749581025E-01-.429010347E-04    3
 .103686234E-07-.655858987E-12-.298390440E+05 .503037294E+02                   4
CYC6H10-O-13            C   6H  10O   1     G    300.00   4000.00 1384.00      1
 .209040427E+02 .249694592E-01-.887525958E-05 .141404459E-08-.835397954E-13    2
-.281106427E+05-.100684615E+03-.120242065E+02 .974927920E-01-.669797836E-04    3
 .211938876E-07-.242310206E-11-.164176421E+05 .774198780E+02                   4
CYC6-OQOOH-3            C   6H  10O   3     G    300.00   4000.00 1421.00      1
 .152391000E+02 .293351956E-01-.936919554E-05 .138764303E-08-.778701917E-13    2
-.379802009E+05-.696293762E+02-.808436864E+01 .898617293E-01-.693837670E-04    3
 .282474384E-07-.463250100E-11-.306468981E+05 .532148412E+02                   4
CYC6-OQOOH-4            C   6H  10O   3     G    300.00   4000.00 1421.00      1
 .152391000E+02 .293351956E-01-.936919554E-05 .138764303E-08-.778701917E-13    2
-.379802009E+05-.703238906E+02-.808436864E+01 .898617293E-01-.693837670E-04    3
 .282474384E-07-.463250100E-11-.306468981E+05 .525203269E+02                   4
ALDEST                  C   6H  10O   3     G    300.00   4000.00 1384.00      1
 .212949599E+02 .266487791E-01-.898035403E-05 .137511216E-08-.789865729E-13    2
-.762788357E+05-.785214726E+02 .521237801E+01 .613142880E-01-.373337900E-04    3
 .119679719E-07-.162337383E-11-.703135588E+05 .903341827E+01                   4
CYC6-OQOOH-2            C   6H  10O   3     G    300.00   4000.00 1416.00      1
 .160913887E+02 .291196520E-01-.940602358E-05 .140488615E-08-.793370497E-13    2
-.378857796E+05-.754185099E+02-.107476916E+02 .986835275E-01-.783513685E-04    3
 .322824282E-07-.532533650E-11-.294335398E+05 .659825481E+02                   4
C6H10O5                 C   6H  10O   5     G    300.00   4000.00 1000.00      1
 .279850422E+02 .264166682E-01-.913640739E-05 .142923991E-08-.833656585E-13    2
-.114313686E+06-.117754445E+03-.781241700E+01 .125424511E+00-.116271866E-03    3
 .544734561E-07-.100746170E-10-.103428291E+06 .690300863E+02                   4
CYC6H12                 C   6H  12          G    300.00   4000.00 1373.00      1
 .190852614E+02 .283866516E-01-.999547753E-05 .158256182E-08-.930877430E-13    2
-.260770569E+05-.880292959E+02-.782903355E+01 .809375102E-01-.439655186E-04    3
 .871887784E-08-.486950162E-15-.157787533E+05 .600472718E+02                   4
NC6H12                  C   6H  12          G    300.00   4000.00 1000.00      1
 .186637886E+02 .209714510E-01-.310828090E-05-.686516180E-09 .160236080E-12    2
-.135910200E+05-.708905467E+02 .196862030E+01 .476562310E-01 .660153730E-05    3
-.371481730E-07 .169224630E-10-.771187890E+04 .208592300E+02                   4
ETBE                    C   6H  14O   1     G    300.00   4000.00 1000.00      1
 .107600227E+02 .484809450E-01-.204693300E-04 .391707780E-08-.279248340E-12    2
-.456695052E+05-.288336460E+02-.321171820E+01 .924083860E-01-.712212230E-04    3
 .295255040E-07-.509148160E-11-.421838470E+05 .417951430E+02                   4
DIPE                    C   6H  14O   1     G    300.00   4000.00 1000.00      1
 .961994133E+01 .527564090E-01-.244349190E-04 .491563770E-08-.360965330E-12    2
-.452985516E+05-.220408754E+02-.207944820E+01 .869029220E-01-.602649600E-04    3
 .209337360E-07-.299614610E-11-.422065600E+05 .378635810E+02                   4
TAME                    C   6H  14O   1     G    300.00   4000.00 1000.00      1
 .102413361E+02 .494717450E-01-.210657300E-04 .406005360E-08-.291140680E-12    2
-.438310029E+05-.257392482E+02-.184725690E+01 .864624650E-01-.624059780E-04    3
 .241227640E-07-.391573010E-11-.407484470E+05 .356637750E+02                   4
C6H5CHO                 C   7H   6O   1     G    300.00   4000.00 1000.00      1
 .151976148E+02 .229544430E-01-.714039470E-05 .736589790E-09 .000000000E+00    2
-.120582935E+05-.546270656E+02-.328352400E+01 .610821620E-01-.279524170E-04    3
 .190203190E-08 .000000000E+00-.599503400E+04 .449259300E+02                   4
C7H8                    C   7H   8          G    300.00   4000.00 1000.00      1
 .988928700E+01 .312351700E-01-.110466410E-04 .129795100E-08 .000000000E+00    2
 .590756417E+03-.294263546E+02-.469518200E+01 .695108030E-01-.438445020E-04    3
 .104046480E-07 .000000000E+00 .469335500E+04 .464073200E+02                   4
CRESOL                  C   7H   8O   1     G    300.00   4000.00 1000.00      1
 .109411883E+02 .359221340E-01-.155859930E-04 .305336930E-08-.221926260E-12    2
-.211837368E+05-.322120090E+02-.410479790E+01 .823735850E-01-.680002460E-04    3
 .287114670E-07-.487123580E-11-.173767210E+05 .440872850E+02                   4
C6H5OCH3                C   7H   8O   1     G    300.00   4000.00 1393.00      1
 .203938728E+02 .209088165E-01-.722522263E-05 .112997840E-08-.659097524E-13    2
-.186061425E+05-.862920505E+02-.540888697E+01 .873332441E-01-.739639658E-04    3
 .320208039E-07-.556946955E-11-.102821510E+05 .500696056E+02                   4
C6H5CH2OH               C   7H   8O   1     G    300.00   4000.00 1000.00      1
 .988928700E+01 .312351700E-01-.110466410E-04 .129795100E-08 .000000000E+00    2
-.176276686E+05-.230348046E+02-.469518200E+01 .695108030E-01-.438445020E-04    3
 .104046480E-07 .000000000E+00-.135250700E+05 .527988700E+02                   4
CH3CH3-C5H6             C   7H  12          G    300.00   4000.00 1000.00      1
 .140192352E+02 .351774100E-01-.121769020E-04 .195853870E-08-.120886390E-12    2
-.562170122E+04-.461295916E+02 .191804150E+01 .620151830E-01-.182958650E-04    3
-.181326460E-07 .113526820E-10-.217165720E+04 .175128710E+02                   4
MCYC6-OQOOH             C   7H  12O   3     G    300.00   4000.00 1380.00      1
 .281047951E+02 .298656134E-01-.103750111E-04 .162883933E-08-.952775107E-13    2
-.587524861E+05-.124642473E+03-.502703972E+01 .104102110E+00-.722526077E-04    3
 .243793077E-07-.320129183E-11-.470307327E+05 .542550536E+02                   4
NC7H14                  C   7H  14          G    300.00   4000.00 1390.00      1
 .206190401E+02 .314852991E-01-.107162057E-04 .165827662E-08-.959911785E-13    2
-.196710875E+05-.822507478E+02-.116533279E+01 .790439806E-01-.496101666E-04    3
 .158569009E-07-.205346433E-11-.117362359E+05 .359871070E+02                   4
MCYC6                   C   7H  14          G    300.00   4000.00 1381.00      1
 .220211359E+02 .332076617E-01-.115857900E-04 .182324838E-08-.106797390E-12    2
-.311719553E+05-.103211614E+03-.890848850E+01 .969226774E-01-.576085500E-04    3
 .148743771E-07-.111357720E-11-.196669630E+05 .657804644E+02                   4
NC7H14O                 C   7H  14O   1     G    300.00   4000.00 1397.00      1
 .231122557E+02 .333659362E-01-.114966228E-04 .179372703E-08-.104427245E-12    2
-.438636425E+05-.993466782E+02-.767475343E+01 .108451023E+00-.827531084E-04    3
 .330380469E-07-.541492429E-11-.334640974E+05 .649157213E+02                   4
NC7H13OOH               C   7H  14O   2     G    300.00   4000.00 1393.00      1
 .277094420E+02 .348487880E-01-.119777002E-04 .186556340E-08-.108475524E-12    2
-.486083259E+05-.114399507E+03 .629165042E+00 .970053636E-01-.668336695E-04    3
 .241186253E-07-.361669837E-11-.390326607E+05 .315310044E+02                   4
NC7-OQOOH               C   7H  14O   3     G    300.00   4000.00 1387.00      1
 .288332529E+02 .320168096E-01-.111508456E-04 .175226159E-08-.102520451E-12    2
-.622309509E+05-.116187714E+03 .152936692E+01 .958173466E-01-.696688520E-04    3
 .269540382E-07-.438728126E-11-.526003608E+05 .306986714E+02                   4
NC7H16                  C   7H  16          G    300.00   4000.00 1000.00      1
 .205103125E+02 .346389640E-01-.107743740E-04 .160399760E-08-.937017530E-13    2
-.326499224E+05-.807081180E+02-.679531340E+00 .810756760E-01-.423279310E-04    3
 .697965770E-08 .837326950E-12-.256907030E+05 .329815600E+02                   4
NC7H15OOH               C   7H  16O   2     G    300.00   4000.00 1393.00      1
 .277094420E+02 .348487880E-01-.119777002E-04 .186556340E-08-.108475524E-12    2
-.486083259E+05-.114399507E+03 .629165042E+00 .970053636E-01-.668336695E-04    3
 .241186253E-07-.361669837E-11-.390326607E+05 .315310044E+02                   4
C8H2                    C   8H   2          G    300.00   4000.00 1000.00      1
 .156802100E+02 .111546100E-01-.372437300E-05 .519789100E-09-.237555000E-13    2
 .108112300E+06-.557143700E+02 .463042700E+01 .393708000E-01-.114803500E-04    3
-.256221400E-07 .167079100E-10 .110828500E+06 .807742500E+00                   4
C6H5C2H                 C   8H   6          G    300.00   4000.00 1399.00      1
 .190886756E+02 .170819066E-01-.559393248E-05 .845345947E-09-.482537486E-13    2
 .280711996E+05-.790035627E+02-.377007730E+01 .792380003E-01-.711832819E-04    3
 .324077613E-07-.583009863E-11 .350595597E+05 .405332699E+02                   4
BZFUR                   C   8H   6O   1     G    300.00   4000.00 1000.00      1
 .161267559E+02 .242942790E-01-.882919089E-05 .143722155E-08-.865592465E-13    2
-.574867958E+04-.640564836E+02-.785221476E+00 .396432449E-01 .569751746E-04    3
-.114831806E-06 .519411145E-10 .215748538E+03 .302655928E+02                   4
C6H5C2H3                C   8H   8          G    300.00   4000.00 1000.00      1
 .132118086E+02 .297097690E-01-.100379980E-04 .113030440E-08 .000000000E+00    2
 .112255113E+05-.452965784E+02-.314842000E+01 .733550410E-01-.482478610E-04    3
 .120551240E-07 .000000000E+00 .157685200E+05 .395339300E+02                   4
XYLENE                  C   8H  10          G    300.00   4000.00 1000.00      1
 .104572604E+02 .403200160E-01-.145441770E-04 .173870560E-08 .000000000E+00    2
-.392485555E+04-.316838798E+02-.365621300E+01 .742185790E-01-.400008720E-04    3
 .741031100E-08 .000000000E+00 .307000000E+03 .427477900E+02                   4
C6H5C2H5                C   8H  10          G    300.00   4000.00 1000.00      1
 .123967254E+02 .365194120E-01-.128125900E-04 .149467160E-08 .000000000E+00    2
-.304290347E+04-.409211516E+02-.458801200E+01 .813929890E-01-.516055260E-04    3
 .123987680E-07 .000000000E+00 .171000000E+04 .472934500E+02                   4
C8H10O3                 C   8H  10O   3     G    300.00   4000.00 1398.00      1
 .397849303E+02 .299091586E-01-.998077835E-05 .152593734E-08-.876494369E-13    2
-.745243570E+05-.176764109E+03-.309175183E+01 .150401311E+00-.141589395E-03    3
 .669336732E-07-.124095424E-10-.617648649E+05 .461394338E+02                   4
UME7                    C   8H  14O   2     G    300.00   4000.00 1386.00      1
 .274195251E+02 .331653074E-01-.112369879E-04 .173174767E-08-.999867016E-13    2
-.597230517E+05-.112624254E+03 .202528941E+01 .898844344E-01-.593620598E-04    3
 .203016355E-07-.286718129E-11-.505953610E+05 .247655861E+02                   4
IC8H16                  C   8H  16          G    300.00   4000.00 1000.00      1
 .159403331E+02 .467083530E-01-.162445520E-04 .262105430E-08-.162114790E-12    2
-.212288474E+05-.575000710E+02-.188446240E+01 .875446570E-01-.337527930E-04    3
-.140196880E-07 .109753600E-10-.160534330E+05 .363096160E+02                   4
IC8H16O                 C   8H  16O   1     G    300.00   4000.00 1400.00      1
 .286870453E+02 .350973257E-01-.120318626E-04 .187165307E-08-.108763411E-12    2
-.489758985E+05-.130519447E+03-.811336944E+01 .120858100E+00-.869108786E-04    3
 .308943900E-07-.431018679E-11-.363657206E+05 .668763983E+02                   4
IC8-OQOOH               C   8H  16O   3     G    300.00   4000.00 1395.00      1
 .329665839E+02 .352889373E-01-.121856584E-04 .190423031E-08-.110989507E-12    2
-.686224367E+05-.138776314E+03 .233137835E+00 .110643301E+00-.779138892E-04    3
 .277663606E-07-.398875833E-11-.571903320E+05 .373387625E+02                   4
IC8H18                  C   8H  18          G    300.00   4000.00 1000.00      1
 .175409498E+02 .499242880E-01-.172020170E-04 .275518900E-08-.169419330E-12    2
-.363533756E+05-.670046390E+02-.203218650E+01 .946845260E-01-.357433050E-04    3
-.165946760E-07 .125346320E-10-.306832730E+05 .359861450E+02                   4
INDENE                  C   9H   8          G    300.00   4000.00 1000.00      1
 .129942100E+02 .345035980E-01-.119473340E-04 .137705200E-08 .000000000E+00    2
 .128398488E+05-.468095535E+02-.565650900E+01 .835992990E-01-.541865810E-04    3
 .131713170E-07 .000000000E+00 .180739000E+05 .501175500E+02                   4
C9H10O2                 C   9H  10O   2     G    300.00   4000.00 1400.00      1
 .279893805E+02 .257305292E-01-.858901356E-05 .131357222E-08-.754726372E-13    2
-.378460988E+05-.119703580E+03-.219761532E+01 .995964750E-01-.769418656E-04    3
 .296736479E-07-.451992280E-11-.279092089E+05 .408797910E+02                   4
TMBENZ                  C   9H  12          G    300.00   4000.00 1383.00      1
 .215885246E+02 .321229102E-01-.110727239E-04 .172825742E-08-.100649304E-12    2
-.136169019E+05-.914142733E+02-.173308850E+01 .786049041E-01-.431048197E-04    3
 .100745302E-07-.585489308E-12-.471446607E+04 .366811038E+02                   4
NPBENZ                  C   9H  12          G    300.00   4000.00 1395.00      1
 .234758956E+02 .300348225E-01-.102493106E-04 .158931255E-08-.921475616E-13    2
-.109980792E+05-.102092892E+03-.597461242E+01 .101439137E+00-.768408376E-04    3
 .299742828E-07-.474668103E-11-.108882285E+04 .550543799E+02                   4
C7H15COCHO              C   9H  16O   2     G    300.00   4000.00 1387.00      1
 .303225194E+02 .381334789E-01-.128450948E-04 .197085647E-08-.113456990E-12    2
-.668175594E+05-.126355483E+03-.229351926E+00 .108754598E+00-.755330139E-04    3
 .275093508E-07-.415197146E-11-.560981532E+05 .380532571E+02                   4
C10H8                   C  10H   8          G    300.00   4000.00 1401.00      1
 .234023214E+02 .242434427E-01-.836282016E-05 .130620111E-08-.761153748E-13    2
 .651941329E+04-.107433208E+03-.883645988E+01 .109300567E+00-.955200914E-04    3
 .421647669E-07-.739851710E-11 .166533366E+05 .621064766E+02                   4
C10H7OH                 C  10H   8O   1     G    300.00   4000.00 1394.00      1
 .262017858E+02 .245473904E-01-.859268465E-05 .135522543E-08-.795056830E-13    2
-.158010339E+05-.119344614E+03-.322687986E+01 .931430619E-01-.687932451E-04    3
 .249753868E-07-.357353464E-11-.568766282E+04 .385570421E+02                   4
C10H10                  C  10H  10          G    300.00   4000.00 2043.00      1
 .196465049E+02 .362867673E-01-.135117921E-04 .222712581E-08-.134868100E-12    2
 .466515480E+04-.883925826E+02-.975555457E+01 .989343734E-01-.593843991E-04    3
 .154882804E-07-.129445409E-11 .148791325E+05 .708155586E+02                   4
TETRALIN                C  10H  12          G    300.00   4000.00 1393.00      1
 .259510150E+02 .311178636E-01-.105072610E-04 .161945272E-08-.935513420E-13    2
-.106963510E+05-.121999608E+03-.103201470E+02 .118533935E+00-.903074920E-04    3
 .343768814E-07-.519161790E-11 .142964373E+04 .715127353E+02                   4
DCYC5                   C  10H  16          G    300.00   4000.00 1396.00      1
 .273482865E+02 .461538793E-01-.158755646E-04 .247442795E-08-.143965250E-12    2
-.380245063E+05-.136978542E+03-.149885463E+02 .144180968E+00-.101905712E-03    3
 .365256640E-07-.527588038E-11-.233132452E+05 .905738933E+02                   4
KHDECA                  C  10H  16O   3     G    300.00   4000.00 1421.00      1
 .152391000E+02 .293351956E-01-.936919554E-05 .138764303E-08-.778701917E-13    2
-.379802009E+05-.703238906E+02-.808436864E+01 .898617293E-01-.693837670E-04    3
 .282474384E-07-.463250100E-11-.306468981E+05 .525203269E+02                   4
DECALIN                 C  10H  18          G    300.00   4000.00 1396.00      1
 .273482865E+02 .461538793E-01-.158755646E-04 .247442795E-08-.143965250E-12    2
-.380245063E+05-.136978542E+03-.149885463E+02 .144180968E+00-.101905712E-03    3
 .365256640E-07-.527588038E-11-.233132452E+05 .905738933E+02                   4
ODECAL                  C  10H  18          G    300.00   4000.00 1383.00      1
 .304308606E+02 .423969327E-01-.145305017E-04 .226051483E-08-.131385276E-12    2
-.274622725E+05-.143201137E+03-.921337866E+01 .127293330E+00-.797537373E-04    3
 .229874961E-07-.227548927E-11-.131010829E+05 .721555536E+02                   4
NC10H20                 C  10H  20          G    300.00   4000.00 1390.00      1
 .306417045E+02 .444757412E-01-.152579717E-04 .237363570E-08-.137907421E-12    2
-.321647483E+05-.129750528E+03-.253770965E+01 .118319727E+00-.776112696E-04    3
 .262647573E-07-.366153318E-11-.202029921E+05 .498650630E+02                   4
NC20MOOH                C  10H  20O   2     G    300.00   4000.00 1393.00      1
 .277094420E+02 .348487880E-01-.119777002E-04 .186556340E-08-.108475524E-12    2
-.486083259E+05-.114399507E+03 .629165042E+00 .970053636E-01-.668336695E-04    3
 .241186253E-07-.361669837E-11-.390326607E+05 .315310044E+02                   4
NC10-OQOOH              C  10H  20O   3     G    300.00   4000.00 1390.00      1
 .373427699E+02 .457774433E-01-.156578702E-04 .243101177E-08-.141046271E-12    2
-.740262240E+05-.156527917E+03 .209018845E+01 .128739739E+00-.918467610E-04    3
 .350282382E-07-.560696315E-11-.617151278E+05 .328016208E+02                   4
NC10H22                 C  10H  22          G    300.00   4000.00 1391.00      1
 .319882239E+02 .477244922E-01-.162276391E-04 .250963259E-08-.145215772E-12    2
-.466392840E+05-.137615344E+03-.208416969E+01 .122535012E+00-.776815739E-04    3
 .249834877E-07-.323548038E-11-.343021863E+05 .471147911E+02                   4
C10H7CHO                C  11H   8O   1     G    300.00   4000.00 1391.00      1
 .276532029E+02 .258287942E-01-.902879433E-05 .142281038E-08-.834251834E-13    2
-.106453206E+05-.124981465E+03-.108527081E+01 .881681978E-01-.575973932E-04    3
 .170999043E-07-.173813923E-11-.356369995E+03 .307785222E+02                   4
C10H7CH3                C  11H  10          G    300.00   4000.00 1394.00      1
 .269623579E+02 .288172394E-01-.100254209E-04 .157466721E-08-.921126923E-13    2
 .586670370E+03-.125206708E+03-.798962224E+01 .117448428E+00-.976360478E-04    3
 .414932114E-07-.710609396E-11 .120022223E+05 .599922187E+02                   4
CH3C10H6OH              C  11H  10O   1     G    300.00   4000.00 1392.00      1
 .281549167E+02 .299236572E-01-.104056239E-04 .163381420E-08-.955470229E-13    2
-.208064399E+05-.126965793E+03-.171335238E+01 .970093442E-01-.665430499E-04    3
 .223717851E-07-.293871610E-11-.102462828E+05 .342637221E+02                   4
C11H12O4                C  11H  12O   4     G    300.00   4000.00 1398.00      1
 .397849303E+02 .299091586E-01-.998077835E-05 .152593734E-08-.876494369E-13    2
-.745243570E+05-.176764109E+03-.309175183E+01 .150401311E+00-.141589395E-03    3
 .669336732E-07-.124095424E-10-.617648649E+05 .461394338E+02                   4
UME10                   C  11H  20O   2     G    300.00   4000.00 1384.00      1
 .374112533E+02 .458948435E-01-.156057696E-04 .241315080E-08-.139673864E-12    2
-.736971925E+05-.162545741E+03 .937241013E+00 .126885097E+00-.836053178E-04    3
 .282312118E-07-.390359926E-11-.605539595E+05 .349335674E+02                   4
ETEROMD                 C  11H  20O   3     G    300.00   4000.00 1386.00      1
 .418053606E+02 .443798286E-01-.151698489E-04 .235874245E-08-.137104681E-12    2
-.896960798E+05-.186388223E+03-.869108022E+00 .143689897E+00-.103700029E-03    3
 .384483018E-07-.582555005E-11-.748416098E+05 .429341731E+02                   4
MDKETO                  C  11H  20O   5     G    300.00   4000.00 1391.00      1
 .435827467E+02 .471875465E-01-.155121189E-04 .235632808E-08-.134947249E-12    2
-.114156459E+06-.184940808E+03 .336575533E+01 .147442203E+00-.113482823E-03    3
 .468018272E-07-.796034235E-11-.100759720E+06 .289177372E+02                   4
MD                      C  11H  22O   2     G    300.00   4000.00 1382.00      1
 .393230373E+02 .488368389E-01-.166923510E-04 .259065840E-08-.150309877E-12    2
-.885441006E+05-.173932688E+03 .176901386E+01 .129360919E+00-.808243357E-04    3
 .251676921E-07-.312062272E-11-.747104475E+05 .304352079E+02                   4
C12H8                   C  12H   8          G    300.00   4000.00 1000.00      1
 .213682716E+02 .324830670E-01-.101214580E-04 .104613640E-08 .000000000E+00    2
 .210494631E+05-.924787980E+02-.672892800E+01 .106967800E+00-.747993040E-04    3
 .193364490E-07 .000000000E+00 .288910000E+05 .533672000E+02                   4
DIBZFUR                 C  12H   8O   1     G    300.00   4000.00 1000.00      1
 .238928699E+02 .342239370E-01-.125916314E-04 .206592304E-08-.125089220E-12    2
-.481449779E+04-.107327684E+03-.194754604E+01 .663215475E-01 .555418713E-04    3
-.135401425E-06 .629515620E-10 .401745217E+04 .350605098E+02                   4
BIPHENYL                C  12H  10          G    300.00   4000.00 1000.00      1
 .214890352E+02 .375797860E-01-.121080230E-04 .129882780E-08 .000000000E+00    2
 .115420788E+05-.916763235E+02-.783196500E+01 .114327200E+00-.776398370E-04    3
 .194042280E-07 .000000000E+00 .198069600E+05 .608493300E+02                   4
DIFENET                 C  12H  10O   1     G    300.00   4000.00 1000.00      1
 .283319364E+02 .317670352E-01-.107447484E-04 .165690065E-08-.957158914E-13    2
-.789446240E+04-.127230446E+03-.865410063E+01 .124988347E+00-.100933530E-03    3
 .413234204E-07-.675938299E-11 .409381103E+04 .686981333E+02                   4
C12H18                  C  12H  18          G    300.00   4000.00 1000.00      1
 .938665800E+02 .198595000E-01-.295692400E-05 .245328200E-09-.917006600E-14    2
-.897187500E+05-.457207000E+03 .374918500E+01 .185852000E+00-.868236800E-04    3
 .615957800E-08 .205893500E-11-.565341800E+05 .387544400E+02                   4
C12H22                  C  12H  22          G    300.00   4000.00 1392.00      1
 .362943970E+02 .488870789E-01-.165740715E-04 .255852468E-08-.147868438E-12    2
-.229987583E+05-.159907963E+03-.329755440E+01 .140713318E+00-.978288195E-04    3
 .352594898E-07-.520523450E-11-.920475977E+04 .529246931E+02                   4
NC12-OQOOH              C  12H  24O   3     G    300.00   4000.00 1678.00      1
 .447068212E+02 .522272795E-01-.195350799E-04 .322923457E-08-.195935332E-12    2
-.818914807E+05-.192299360E+03 .877388676E+01 .119113497E+00-.561329021E-04    3
 .677643630E-08 .106366869E-11-.685051188E+05 .572134782E+01                   4
NC12H26                 C  12H  26          G    300.00   4000.00 1391.00      1
 .385099212E+02 .563550048E-01-.191493200E-04 .296024862E-08-.171244150E-12    2
-.548849270E+05-.169785166E+03-.262181594E+01 .147237711E+00-.943970271E-04    3
 .307441268E-07-.403602230E-11-.400654253E+05 .529882396E+02                   4
FLUORENE                C  13H  10          G    300.00   4000.00 1000.00      1
 .231612871E+02 .392128530E-01-.125431510E-04 .133503890E-08 .000000000E+00    2
 .123102892E+05-.103717257E+03-.112092800E+02 .129847800E+00-.907013380E-04    3
 .232288460E-07 .000000000E+00 .219426600E+05 .748524200E+02                   4
C6H5CH2C6H5             C  13H  12          G    300.00   4000.00 1000.00      1
 .185418955E+02 .513343070E-01-.178726910E-04 .207043850E-08 .000000000E+00    2
 .668552054E+04-.690121392E+02-.940899900E+01 .125451300E+00-.822539730E-04    3
 .202856220E-07 .000000000E+00 .144845500E+05 .760677200E+02                   4
ALDINS                  C  13H  20O   1     G    300.00   4000.00 1000.00      1
 .938665800E+02 .198595000E-01-.295692400E-05 .245328200E-09-.917006600E-14    2
-.897187500E+05-.457207000E+03 .374918500E+01 .185852000E+00-.868236800E-04    3
 .615957800E-08 .205893500E-11-.565341800E+05 .387544400E+02                   4
U2ME12                  C  13H  22O   2     G    300.00   4000.00 1391.00      1
 .422353117E+02 .524987045E-01-.181261023E-04 .283174793E-08-.165001495E-12    2
-.676968189E+05-.186270028E+03 .679798314E-01 .152530074E+00-.111376081E-03    3
 .435663556E-07-.715842617E-11-.529996239E+05 .399987338E+02                   4
C14H10                  C  14H  10          G    300.00   4000.00 1000.00      1
 .255171870E+02 .393727940E-01-.123155080E-04 .127852800E-08 .000000000E+00    2
 .131224037E+05-.115618425E+03-.909474100E+01 .131333800E+00-.924017290E-04    3
 .240156710E-07 .000000000E+00 .227649500E+05 .639753600E+02                   4
C6H5C2H4C6H5            C  14H  14          G    300.00   4000.00 1000.00      1
 .183724857E+02 .606470630E-01-.215506390E-04 .254284330E-08 .000000000E+00    2
 .518516081E+04-.659251182E+02-.814781700E+01 .130620600E+00-.819367560E-04    3
 .194757260E-07 .000000000E+00 .126141800E+05 .718458700E+02                   4
C16H10                  C  16H  10          G    300.00   4000.00 1000.00      1
 .290747022E+02 .412337670E-01-.126077060E-04 .127453580E-08 .000000000E+00    2
 .141687238E+05-.136431347E+03-.106811200E+02 .146535400E+00-.103943520E-03    3
 .270645390E-07 .000000000E+00 .252715000E+05 .699617500E+02                   4
NC16-OQOOH              C  16H  32O   3     G    300.00   4000.00 1854.00      1
 .488264318E+02 .825357366E-01-.292747409E-04 .467245514E-08-.276718037E-12    2
-.942845289E+05-.205583924E+03 .138386904E+01 .198379105E+00-.134722947E-03    3
 .475955890E-07-.691333208E-11-.791319641E+05 .463051187E+02                   4
IC16-OQOOH              C  16H  32O   3     G    300.00   4000.00 1397.00      1
 .620188250E+02 .682375774E-01-.235322180E-04 .367416933E-08-.214025539E-12    2
-.107194396E+06-.296402060E+03-.700111687E+01 .236135134E+00-.181200158E-03    3
 .715715364E-07-.114883341E-10-.839739066E+05 .717765001E+02                   4
NC16H34                 C  16H  34          G    300.00   4000.00 1391.00      1
 .515593854E+02 .736064257E-01-.249888737E-04 .386085377E-08-.223263662E-12    2
-.713781425E+05-.234158439E+03-.369111950E+01 .196612966E+00-.127777824E-03    3
 .422323349E-07-.562967041E-11-.515927302E+05 .647080513E+02                   4
IC16H34                 C  16H  34          G    300.00   4000.00 1400.00      1
 .565856523E+02 .692869560E-01-.234931111E-04 .362720220E-08-.209665225E-12    2
-.820366778E+05-.276851694E+03-.107545408E+02 .233995831E+00-.178076331E-03    3
 .696956034E-07-.110282035E-10-.595981394E+05 .818346760E+02                   4
UME16                   C  17H  32O   2     G    300.00   4000.00 1000.00      1
 .333606142E+02 .106719124E+00-.429500189E-04 .790457654E-08-.546125152E-12    2
-.868236054E+05-.126816968E+03 .114310960E+02 .102101194E+00 .102480878E-03    3
-.181385357E-06 .698603588E-10-.778209017E+05 .206428096E+01                   4
ETEROMPA                C  17H  32O   3     G    300.00   4000.00 1000.00      1
 .406345250E+02 .963702350E-01-.332815250E-04 .536978820E-08-.333546480E-12    2
-.105022900E+06-.161181400E+03-.374618910E+01 .216936450E+00-.134184780E-03    3
 .217036750E-07 .800116570E-11-.930412810E+05 .677468110E+02                   4
MPA                     C  17H  34O   2     G    300.00   4000.00 1000.00      1
 .355305296E+02 .109746228E+00-.440981772E-04 .810571172E-08-.559469785E-12    2
-.102923616E+06-.145292419E+03 .117629996E+02 .108027697E+00 .103662595E-03    3
-.187190120E-06 .724616510E-10-.933306777E+05-.643066315E+01                   4
KHMLIN1                 C  19H  30O   5     G    300.00   4000.00 1843.00      1
 .597680898E+02 .832144998E-01-.302817533E-04 .491632066E-08-.294624551E-12    2
-.961002787E+05-.258440317E+03-.347354324E+01 .238348931E+00-.171810701E-03    3
 .624560833E-07-.914836595E-11-.760003616E+05 .770024622E+02                   4
MLIN1                   C  19H  32O   2     G    300.00   4000.00 1834.00      1
 .520202170E+02 .871284776E-01-.313984409E-04 .506450961E-08-.302130761E-12    2
-.727531890E+05-.226713941E+03-.298592567E+01 .218746556E+00-.148096154E-03    3
 .511216154E-07-.719451974E-11-.549290521E+05 .662774857E+02                   4
MLINO                   C  19H  34O   2     G    300.00   4000.00 1833.00      1
 .524257963E+02 .910351615E-01-.326514183E-04 .524998946E-08-.312507814E-12    2
-.869039436E+05-.227879204E+03-.158761924E+01 .219526542E+00-.145761172E-03    3
 .495347572E-07-.688636525E-11-.693288124E+05 .600962817E+02                   4
MEOLE                   C  19H  36O   2     G    300.00   4000.00 1831.00      1
 .528856562E+02 .948572658E-01-.338668063E-04 .542873444E-08-.322458135E-12    2
-.101075125E+06-.229348639E+03-.267573662E+00 .220639742E+00-.143861659E-03    3
 .481699649E-07-.661786902E-11-.837166223E+05 .542791001E+02                   4
MSTEAKETO               C  19H  36O   5     G    300.00   4000.00 1857.00      1
 .628573476E+02 .927885184E-01-.331648431E-04 .532086973E-08-.316267196E-12    2
-.142644021E+06-.277684268E+03-.711176329E+00 .251338095E+00-.180571731E-03    3
 .664483461E-07-.990089173E-11-.122716422E+06 .585265768E+02                   4
MSTEA                   C  19H  38O   2     G    300.00   4000.00 1000.00      1
 .418174710E+02 .117959830E+00-.465265590E-04 .845319460E-08-.579171090E-12    2
-.110862900E+06-.175601040E+03 .114771030E+02 .131225240E+00 .898738730E-04    3
-.183685190E-06 .722337400E-10-.991500330E+05-.163992920E+01                   4
BIN1B                   C  20H  10          G    300.00   4000.00 1000.00      1
-.570256700E+01 .143432300E+00-.880724700E-04 .276799200E-07-.352289900E-11    2
 .277808900E+05 .434481200E+02-.570256700E+01 .143432300E+00-.880724700E-04    3
 .276799200E-07-.352289900E-11 .277808900E+05 .434481200E+02                   4
BIN1A                   C  20H  16          G    300.00   4000.00 1000.00      1
-.324173600E+01 .158222900E+00-.946183500E-04 .281843100E-07-.356131000E-11    2
 .217869900E+05 .300825300E+02-.324173600E+01 .158222900E+00-.946183500E-04    3
 .281843100E-07-.356131000E-11 .217869900E+05 .300825300E+02                   4
N                       N   1               G    300.00   4000.00 1000.00      1
 .245026778E+01 .106614600E-03-.746533710E-07 .187965200E-10-.102598400E-14    2
 .561160257E+05 .444874779E+01 .250307100E+01-.218001810E-04 .542052910E-07    3
-.564755990E-10 .209990390E-13 .560988900E+05 .416756600E+01                   4
O                       O   1               G    300.00   4000.00 1000.00      1
 .254205876E+01-.275506100E-04-.310280290E-08 .455106700E-11-.436805100E-15    2
 .292307989E+05 .492030884E+01 .294642800E+01-.163816600E-02 .242103100E-05    3
-.160284300E-08 .389069610E-12 .291476400E+05 .296399500E+01                   4
NO3                     O   3N   1          G    300.00   4000.00 1000.00      1
 .712030587E+01 .324622800E-02-.143161340E-05 .279705300E-09-.201300700E-13    2
 .586448126E+04-.121372920E+02 .122107630E+01 .187879700E-01-.134432120E-04    3
 .127460130E-08 .135406010E-11 .747314400E+04 .184020200E+02                   4
H                       H   1               G    300.00   4000.00 1000.00      1
 .250000000E+01 .000000000E+00 .000000000E+00 .000000000E+00 .000000000E+00    2
 .254716200E+05-.460117600E+00 .250000000E+01 .000000000E+00 .000000000E+00    3
 .000000000E+00 .000000000E+00 .254716200E+05-.460117600E+00                   4
NH                      H   1N   1          G    300.00   4000.00 1000.00      1
 .276025108E+01 .137534600E-02-.445191400E-06 .769279080E-10-.501759190E-14    2
 .420782748E+05 .585718609E+01 .333975800E+01 .125300900E-02-.349164500E-05    3
 .421881200E-08-.155761800E-11 .418504700E+05 .250718000E+01                   4
NNH                     H   1N   2          G    300.00   4000.00 1000.00      1
 .441534072E+01 .161438800E-02-.163289400E-06-.855984590E-10 .161479110E-13    2
 .278802961E+05 .904297112E+00 .350134400E+01 .205358610E-02 .717040900E-06    3
 .492134780E-09-.967117010E-12 .283334700E+05 .639183800E+01                   4
OH                      H   1O   1          G    300.00   4000.00 1710.00      1
 .285376040E+01 .102994334E-02-.232666477E-06 .193750704E-10-.315759847E-15    2
 .369949720E+04 .578756825E+01 .341896226E+01 .319255801E-03-.308292717E-06    3
 .364407494E-09-.100195479E-12 .345264448E+04 .254433372E+01                   4
HO2                     H   1O   2          G    300.00   4000.00 1000.00      1
 .401721090E+01 .223982013E-02-.633658150E-06 .114246370E-09-.107908535E-13    2
 .111856713E+03 .378510215E+01 .430179801E+01-.474912051E-02 .211582891E-04    3
-.242763894E-07 .929225124E-11 .294808040E+03 .371666245E+01                   4
NH2                     H   2N   1          G    300.00   4000.00 1000.00      1
 .296131091E+01 .293269890E-02-.906360010E-06 .161725700E-09-.120420000E-13    2
 .219197637E+05 .577788090E+01 .343249300E+01 .329953990E-02-.661359990E-05    3
 .859094660E-08-.357204610E-11 .217722700E+05 .309011000E+01                   4
H2NO                    H   2O   1N   1     G    300.00   4000.00 1000.00      1
 .149675000E+01 .889472000E-02-.330837000E-05 .405760000E-09 .000000000E+00    2
 .724825208E+04 .175864616E+02 .267141000E+01 .529823000E-02 .360637000E-06    3
-.841417000E-09 .000000000E+00 .696062900E+04 .116499100E+02                   4
N2H3                    H   3N   2          G    300.00   4000.00 1000.00      1
 .444184100E+01 .721427100E-02-.249568400E-05 .392056500E-09-.229895000E-13    2
 .166422164E+05-.427486304E+00 .317420400E+01 .471590700E-02 .133486700E-04    3
-.191968500E-07 .748756400E-11 .172727000E+05 .755722400E+01                   4
CSOLID                  C   1               G    300.00   4000.00 1000.00      1
 .145569246E+01 .171706380E-02-.697584100E-06 .135283160E-09-.967649050E-14    2
-.695128087E+03-.852568475E+01-.310872070E+00 .440353690E-02 .190394120E-05    3
-.638546970E-08 .298964250E-11-.108650790E+03 .111382950E+01                   4
C                       C   1               G    300.00   4000.00 1000.00      1
 .249266888E+01 .479889284E-04-.724335020E-07 .374291029E-10-.487277893E-14    2
 .854512953E+05 .480150373E+01 .255423955E+01-.321537724E-03 .733792245E-06    3
-.732234889E-09 .266521446E-12 .854438832E+05 .453130848E+01                   4
CN                      C   1N   1          G    300.00   4000.00 1000.00      1
 .372011754E+01 .151835110E-03 .198738110E-06-.379837100E-10 .132823000E-14    2
 .511162563E+05 .288861031E+01 .366320400E+01-.115652890E-02 .216340890E-05    3
 .185420800E-09-.821469520E-12 .512811700E+05 .373901500E+01                   4
NCO                     C   1O   1N   1     G    300.00   4000.00 1000.00      1
 .501204558E+01 .262677300E-02-.110824310E-05 .209385990E-09-.146034700E-13    2
 .173718555E+05-.183007911E+01 .283032000E+01 .887149010E-02-.894563620E-05    3
 .587691810E-08-.190773400E-11 .180054300E+05 .949883200E+01                   4
CH                      C   1H   1          G    300.00   4000.00 1000.00      1
 .219622115E+01 .234038100E-02-.705820130E-06 .900758220E-10-.385504010E-14    2
 .708672121E+05 .917838138E+01 .320020200E+01 .207287490E-02-.513443090E-05    3
 .573388980E-08-.195553300E-11 .704525700E+05 .333158700E+01                   4
HCO                     C   1H   1O   1     G    300.00   4000.00 1000.00      1
 .355727119E+01 .334557190E-02-.133500600E-05 .247057210E-09-.171385000E-13    2
 .391632208E+04 .555229973E+01 .289832900E+01 .619914620E-02-.962308420E-05    3
 .108982500E-07-.457488520E-11 .415992100E+04 .898361500E+01                   4
HCO3                    C   1H   1O   3     G    300.00   4000.00 1368.00      1
 .724073447E+01 .463312951E-02-.163693995E-05 .259706693E-09-.152964699E-13    2
-.187027386E+05-.649534993E+01 .396059309E+01 .106002279E-01-.525713351E-05    3
 .101716726E-08-.287487602E-13-.173599383E+05 .117807483E+02                   4
CH2S                    C   1H   2          G    300.00   4000.00 1000.00      1
 .355288641E+01 .206678800E-02-.191411600E-06-.110467300E-09 .202134890E-13    2
 .498497521E+05 .168658499E+01 .397126500E+01-.169908800E-03 .102536900E-05    3
 .249254990E-08-.198126610E-11 .498936700E+05 .575320760E-01                   4
CH2                     C   1H   2          G    300.00   4000.00 1000.00      1
 .363640757E+01 .193305600E-02-.168701600E-06-.100989900E-09 .180825510E-13    2
 .453413341E+05 .215656196E+01 .376223700E+01 .115981900E-02 .248958490E-06    3
 .880083620E-09-.733243490E-12 .453679000E+05 .171257700E+01                   4
H2CN                    C   1H   2N   1     G    300.00   4000.00 1000.00      1
 .520970151E+01 .296929110E-02-.285558910E-06-.163555000E-09 .304325890E-13    2
 .276771105E+05-.444446452E+01 .285166100E+01 .569523310E-02 .107114000E-05    3
-.162261200E-08-.235110810E-12 .286378200E+05 .899274900E+01                   4
CH3                     C   1H   3          G    300.00   4000.00 1000.00      1
 .284405718E+01 .613797410E-02-.223034500E-05 .378516110E-09-.245215900E-13    2
 .164378004E+05 .545265727E+01 .243044200E+01 .111241000E-01-.168022000E-04    3
 .162182910E-07-.586495220E-11 .164237800E+05 .678979400E+01                   4
CH3O                    C   1H   3O   1     G    300.00   4000.00 1000.00      1
 .377081447E+01 .787149740E-02-.265638390E-05 .394443090E-09-.211261600E-13    2
 .127818951E+03 .292947482E+01 .210620400E+01 .721659510E-02 .533847200E-05    3
-.737763630E-08 .207561010E-11 .978601200E+03 .131521800E+02                   4
CH2OH                   C   1H   3O   1     G    300.00   4000.00 1000.00      1
 .632751914E+01 .360827010E-02-.320154700E-06-.193875000E-09 .350970410E-13    2
-.447450931E+04-.832935988E+01 .286262800E+01 .100152700E-01-.528543520E-06    3
-.513853890E-08 .224604100E-11-.334967800E+04 .103979400E+02                   4
CH3OO                   C   1H   3O   2     G    300.00   4000.00 1385.00      1
 .595784570E+01 .790728626E-02-.268246234E-05 .413891337E-09-.239007330E-13    2
-.378178515E+03-.353671121E+01 .426146906E+01 .100873599E-01-.321506184E-05    3
 .209409267E-09 .418339103E-13 .473129653E+03 .634599067E+01                   4
C2H                     C   2H   1          G    300.00   4000.00 1000.00      1
 .316780603E+01 .475221900E-02-.183787070E-05 .304190250E-09-.177232770E-13    2
 .671210651E+05 .663589763E+01 .288965730E+01 .134099610E-01-.284769500E-04    3
 .294791040E-07-.109331510E-10 .668393930E+05 .622296430E+01                   4
HCCO                    C   2H   1O   1     G    300.00   4000.00 1000.00      1
 .675807437E+01 .200040010E-02-.202760700E-06-.104113200E-09 .196516400E-13    2
 .190151261E+05-.907126528E+01 .504796600E+01 .445347790E-02 .226828210E-06    3
-.148209400E-08 .225074100E-12 .196589100E+05 .481843900E+00                   4
CH2CN                   C   2H   2N   1     G    300.00   4000.00 1000.00      1
 .460581482E+01 .944851600E-02-.471163290E-05 .113899570E-08-.108289420E-12    2
 .291714861E+05 .100843943E+01 .252967240E+01 .181141380E-01-.189605750E-04    3
 .119445830E-07-.325441420E-11 .295922930E+05 .109934410E+02                   4
C2H3                    C   2H   3          G    300.00   4000.00 1000.00      1
 .593346697E+01 .401774510E-02-.396673900E-06-.144126700E-09 .237864300E-13    2
 .318543468E+05-.853030497E+01 .245927600E+01 .737147590E-02 .210987200E-05    3
-.132164200E-08-.118478400E-11 .333522500E+05 .115562000E+02                   4
CH3CO                   C   2H   3O   1     G    300.00   4000.00 1000.00      1
 .561230883E+01 .844988600E-02-.285414690E-05 .423837600E-09-.226840300E-13    2
-.518788372E+04-.327515155E+01 .312527800E+01 .977822020E-02 .452144790E-05    3
-.900946160E-08 .319371700E-11-.410850700E+04 .112288500E+02                   4
CH2CHO                  C   2H   3O   1     G    300.00   4000.00 1500.00      1
 .971005743E+01 .385496600E-02-.467782500E-06-.150517900E-09 .294142800E-13    2
-.269248263E+04-.281056408E+02 .280220500E+00 .274031100E-01-.255468300E-04    3
 .130667900E-07-.275042500E-11 .668264800E+03 .223973100E+02                   4
CH3OCO                  C   2H   3O   2     G    300.00   4000.00 1601.00      1
 .973659803E+01 .742432713E-02-.265641779E-05 .425031143E-09-.251824924E-13    2
-.235512450E+05-.237360013E+02 .416215406E+01 .138037511E-01-.308486109E-06    3
-.456430814E-08 .146909632E-11-.209627030E+05 .854235619E+01                   4
CH3CO3                  C   2H   3O   3     G    300.00   4000.00 1000.00      1
 .102188027E+02 .888408630E-02-.222887620E-05 .166265570E-09 .000000000E+00    2
-.256023886E+05-.219354293E+02 .384065500E+01 .218595100E-01-.904528040E-05    3
 .385393800E-09 .000000000E+00-.234946000E+05 .124829900E+02                   4
C2H5                    C   2H   5          G    300.00   4000.00 1000.00      1
 .719047846E+01 .648407680E-02-.642806410E-06-.234787910E-09 .388087690E-13    2
 .106745471E+05-.147808755E+02 .269070100E+01 .871913320E-02 .441983820E-05    3
 .933870310E-09-.392777300E-11 .128704000E+05 .121382000E+02                   4
C2H4OH                  C   2H   5O   1     G    300.00   4000.00 1391.00      1
 .752244726E+01 .110492715E-01-.372576465E-05 .572827397E-09-.330061759E-13    2
-.729337464E+04-.124960750E+02 .117714711E+01 .248115685E-01-.150299503E-04    3
 .479006785E-08-.640994211E-12-.495369043E+04 .220081586E+02                   4
CH3OCH2                 C   2H   5O   1     G    300.00   4000.00 1376.00      1
 .817131769E+01 .110086181E-01-.382352277E-05 .599637202E-09-.350317513E-13    2
-.291606126E+04-.178646468E+02 .291327415E+01 .203364659E-01-.959712342E-05    3
 .207478525E-08-.171343362E-12-.685171134E+03 .116066817E+02                   4
CH3CHOH                 C   2H   5O   1     G    300.00   4000.00 1553.00      1
 .726570301E+01 .109588926E-01-.363662803E-05 .553659830E-09-.317012322E-13    2
-.864371441E+04-.106822851E+02 .183974631E+01 .187789371E-01-.460544253E-05    3
-.213116990E-08 .943772653E-12-.629595195E+04 .201446141E+02                   4
C2H5OO                  C   2H   5O   2     G    300.00   4000.00 1388.00      1
 .951115499E+01 .122676900E-01-.422364452E-05 .658474989E-09-.383095208E-13    2
-.676067578E+04-.223427083E+02 .177950508E+01 .304938087E-01-.216376209E-04    3
 .868906296E-08-.151788464E-11-.399101974E+04 .192919501E+02                   4
C2-QOOH                 C   2H   5O   2     G    300.00   4000.00 1396.00      1
 .116258666E+02 .100826346E-01-.347934362E-05 .543394220E-09-.316569294E-13    2
-.910568267E+03-.318522902E+02 .813237801E+00 .390063400E-01-.340643855E-04    3
 .155066226E-07-.284069840E-11 .250785787E+04 .249684459E+02                   4
DME-OO                  C   2H   5O   3     G    300.00   4000.00 1359.00      1
 .120501213E+02 .123072703E-01-.435221905E-05 .690896352E-09-.407091104E-13    2
-.227977573E+05-.323415629E+02 .515628105E+01 .216783339E-01-.561847228E-05    3
-.192807296E-08 .859447044E-12-.196244836E+05 .725163812E+01                   4
DME-QOOH                C   2H   5O   3     G    300.00   4000.00 1367.00      1
 .140894827E+02 .105710448E-01-.375281006E-05 .597314407E-09-.352604582E-13    2
-.191406716E+05-.429268872E+02 .543520255E+01 .272005914E-01-.150210893E-04    3
 .370396290E-08-.309396378E-12-.157034464E+05 .495012674E+01                   4
C2-OOQOOH               C   2H   5O   4     G    300.00   4000.00 1387.00      1
 .145471032E+02 .123393823E-01-.427259469E-05 .668763337E-09-.390196721E-13    2
-.196338761E+05-.408784236E+02 .590031872E+01 .305658528E-01-.185905950E-04    3
 .567871605E-08-.702799577E-12-.163916571E+05 .633051038E+01                   4
DME-OOQOOH              C   2H   5O   5     G    300.00   4000.00 1382.00      1
 .146274659E+02 .163794767E-01-.563311171E-05 .877481381E-09-.510186598E-13    2
-.370029335E+05-.399555488E+02 .771229157E+01 .301140957E-01-.165996092E-04    3
 .533577253E-08-.842885930E-12-.341808026E+05-.165902348E+01                   4
C3H3                    C   3H   3          G    300.00   4000.00 1000.00      1
 .883104772E+01 .435719410E-02-.410906610E-06-.236872300E-09 .437652000E-13    2
 .384741917E+05-.217791939E+02 .475419900E+01 .110802800E-01 .279332310E-06    3
-.547921220E-08 .194962900E-11 .398888300E+05 .585454700E+00                   4
CH2CHCH2                C   3H   5          G    300.00   4000.00 1000.00      1
 .846871473E+01 .110576240E-01-.329817360E-05 .323385870E-09 .000000000E+00    2
 .160467269E+05-.206696057E+02 .227648600E+01 .198556410E-01 .112384200E-05    3
-.101457600E-07 .344134200E-11 .182949600E+05 .137251500E+02                   4
CH2CCH3                 C   3H   5          G    300.00   4000.00 1000.00      1
 .920976624E+01 .787141170E-02-.772452210E-06-.449735690E-09 .837727170E-13    2
 .285396699E+05-.223237088E+02 .316186300E+01 .151810000E-01 .272265900E-05    3
-.517711210E-08 .543528610E-13 .309554700E+05 .119797300E+02                   4
CHCHCH3                 C   3H   5          G    300.00   4000.00 1000.00      1
 .920976624E+01 .787141170E-02-.772452210E-06-.449735690E-09 .837727170E-13    2
 .285396699E+05-.223237088E+02 .316186300E+01 .151810000E-01 .272265900E-05    3
-.517711210E-08 .543528610E-13 .309554700E+05 .119797300E+02                   4
C2H4CHO                 C   3H   5O   1     G    300.00   4000.00 1683.00      1
 .813285396E+01 .137651720E-01-.486366739E-05 .775334875E-09-.459117207E-13    2
-.292071282E+04-.132464943E+02 .324839539E+01 .209600531E-01-.607665825E-05    3
-.115341896E-08 .627874009E-12-.913395491E+03 .143591941E+02                   4
CH3COCH2                C   3H   5O   1     G    300.00   4000.00 1391.00      1
 .102303674E+02 .116494161E-01-.401005537E-05 .625205246E-09-.363784362E-13    2
-.844376284E+04-.279195044E+02 .180339187E+01 .301407085E-01-.193505552E-04    3
 .638199034E-08-.866103180E-12-.537233261E+04 .178046408E+02                   4
C3H5OO                  C   3H   5O   2     G    300.00   4000.00 1375.00      1
 .120289627E+02 .126220050E-01-.443107280E-05 .699998849E-09-.411059161E-13    2
 .440592543E+04-.346276747E+02 .316765415E+01 .300862111E-01-.169786280E-04    3
 .462955698E-08-.501220245E-12 .789477349E+04 .142601307E+02                   4
IC3H7                   C   3H   7          G    300.00   4000.00 1000.00      1
 .736341098E+01 .171331520E-01-.582028000E-05 .658834320E-09 .000000000E+00    2
 .604684608E+04-.148406654E+02 .171329900E+01 .254261610E-01 .158080800E-05    3
-.182128610E-07 .882771030E-11 .803580600E+04 .162790100E+02                   4
NC3H7                   C   3H   7          G    300.00   4000.00 1000.00      1
 .722715260E+01 .172648710E-01-.588880490E-05 .669183600E-09 .000000000E+00    2
 .782835831E+04-.127978858E+02 .192253600E+01 .247892700E-01 .181024900E-05    3
-.178326490E-07 .858299630E-11 .971328300E+04 .164927100E+02                   4
CH3CH2CH2O              C   3H   7O   1     G    300.00   4000.00 1386.00      1
 .114171877E+02 .153513978E-01-.529698955E-05 .827233821E-09-.481919070E-13    2
-.102618580E+05-.351878119E+02 .408331131E+00 .386748099E-01-.236531335E-04    3
 .722163698E-08-.882900722E-12-.615994143E+04 .248520294E+02                   4
CH2CH2CH2OH             C   3H   7O   1     G    300.00   4000.00 1392.00      1
 .106573810E+02 .155684549E-01-.527663821E-05 .814099260E-09-.470228616E-13    2
-.112728087E+05-.272448749E+02 .975268381E+00 .369225253E-01-.232066980E-04    3
 .768472523E-08-.106762046E-11-.774554528E+04 .252661698E+02                   4
CH2CHOHCH3              C   3H   7O   1     G    300.00   4000.00 1388.00      1
 .110944203E+02 .153549108E-01-.523574640E-05 .810964124E-09-.469665855E-13    2
-.134769536E+05-.307070215E+02 .584672920E+00 .407370189E-01-.294865043E-04    3
 .116950656E-07-.196228356E-11-.984929391E+04 .255429190E+02                   4
CH3CHCH2OH              C   3H   7O   1     G    300.00   4000.00 1674.00      1
 .931287816E+01 .167579212E-01-.575555480E-05 .900584362E-09-.526566836E-13    2
-.119163093E+05-.195564662E+02 .120494302E+01 .330857885E-01-.163893637E-04    3
 .318103918E-08-.684229288E-13-.902896295E+04 .246601603E+02                   4
CH3CH2CHOH              C   3H   7O   1     G    300.00   4000.00 1386.00      1
 .110500439E+02 .152562747E-01-.517257413E-05 .798146428E-09-.461030406E-13    2
-.142779432E+05-.312276095E+02 .149130595E+01 .376502110E-01-.258507542E-04    3
 .978662277E-08-.158835656E-11-.109017244E+05 .201908977E+02                   4
NC3H7O                  C   3H   7O   1     G    300.00   4000.00 1390.00      1
 .107032043E+02 .160908541E-01-.548805425E-05 .850429828E-09-.492755368E-13    2
-.101405419E+05-.313058764E+02-.595838475E+00 .410450833E-01-.263340323E-04    3
 .872638287E-08-.119115039E-11-.604569631E+04 .299328965E+02                   4
CH3COHCH3               C   3H   7O   1     G    300.00   4000.00 1388.00      1
 .115026438E+02 .149881248E-01-.510421075E-05 .789864272E-09-.457135659E-13    2
-.164821894E+05-.347655748E+02 .118802517E+01 .410410262E-01-.314650841E-04    3
 .133514692E-07-.237788249E-11-.130177234E+05 .200655998E+02                   4
NC3H7OO                 C   3H   7O   2     G    300.00   4000.00 1388.00      1
 .127230991E+02 .167336808E-01-.575943184E-05 .897769493E-09-.522275065E-13    2
-.108816595E+05-.381965321E+02 .156301709E+01 .426192697E-01-.296615075E-04    3
 .114187326E-07-.189894471E-11-.688086375E+04 .219842933E+02                   4
IC3H7OO                 C   3H   7O   2     G    300.00   4000.00 1392.00      1
 .132610651E+02 .162501084E-01-.558631798E-05 .870057473E-09-.505849469E-13    2
-.131937089E+05-.421023499E+02 .103495454E+01 .469942369E-01-.366525520E-04    3
 .157084173E-07-.281956117E-11-.906344820E+04 .229566921E+02                   4
IC3-QOOH                C   3H   7O   2     G    300.00   4000.00 1399.00      1
 .155030898E+02 .139802008E-01-.481811216E-05 .751835399E-09-.437743118E-13    2
-.741643030E+04-.523911482E+02-.184042862E+00 .564670638E-01-.501611253E-04    3
 .230526863E-07-.423866481E-11-.252333896E+04 .298354826E+02                   4
NC3-QOOH                C   3H   7O   2     G    300.00   4000.00 1374.00      1
 .146139980E+02 .143723015E-01-.488635144E-05 .756519620E-09-.438364992E-13    2
-.646101457E+04-.457478245E+02 .191005011E+01 .411666833E-01-.251630217E-04    3
 .711856873E-08-.698838732E-12-.179305093E+04 .234514457E+02                   4
IC3-OOQOOH              C   3H   7O   4     G    300.00   4000.00 1391.00      1
 .191234208E+02 .158457151E-01-.552231946E-05 .868162288E-09-.508094203E-13    2
-.255253957E+05-.661419362E+02 .175906535E+01 .624712381E-01-.554930416E-04    3
 .257973727E-07-.483190839E-11-.200009572E+05 .251348546E+02                   4
NC3-OOQOOH              C   3H   7O   4     G    300.00   4000.00 1388.00      1
 .185146106E+02 .164157074E-01-.573085844E-05 .901975314E-09-.528299084E-13    2
-.231819444E+05-.618247164E+02 .254387733E+01 .570847379E-01-.472164204E-04    3
 .208289492E-07-.378162942E-11-.178600410E+05 .229447574E+02                   4
C4H3                    C   4H   3          G    300.00   4000.00 1000.00      1
 .107527376E+02 .538115300E-02-.554963720E-06-.305226590E-09 .576173970E-13    2
 .612141980E+05-.297302533E+02 .415388100E+01 .172628700E-01-.238937390E-06    3
-.101870000E-07 .434050410E-11 .633807200E+05 .603650600E+01                   4
C4H3O                   C   4H   3O   1     G    300.00   4000.00 1000.00      1
 .129455763E+02 .795235476E-02-.280679691E-05 .445205248E-09-.262240810E-13    2
 .175946397E+05-.478819894E+02-.584674088E+01 .620875882E-01-.630010605E-04    3
 .306882361E-07-.575456234E-11 .230253176E+05 .492940922E+02                   4
C4H5                    C   4H   5          G    300.00   4000.00 1000.00      1
 .128659744E+02 .794336940E-02-.862646570E-06-.465563500E-09 .895113110E-13    2
 .378355213E+05-.418250446E+02 .299524000E+01 .228845610E-01 .197547090E-05    3
-.114824500E-07 .319782310E-11 .414221800E+05 .128945400E+02                   4
IC4H7                   C   4H   7          G    300.00   4000.00 1000.00      1
 .616543300E+01 .257842760E-01-.936521250E-05 .112618500E-08 .000000000E+00    2
 .114713700E+05-.676561500E+01 .476952000E+01 .167724920E-01 .213011010E-04    3
-.275874430E-07 .845501100E-11 .126384700E+05 .401309300E+01                   4
SC4H7                   C   4H   7          G    300.00   4000.00 1000.00      1
 .714879043E+01 .219663880E-01-.774471300E-05 .907477370E-09 .000000000E+00    2
 .124589843E+05-.117547735E+02-.442598200E+00 .422160100E-01-.254697900E-04    3
 .597432100E-08 .000000000E+00 .145672100E+05 .276086500E+02                   4
CH2C3H5                 C   4H   7          G    300.00   4000.00 1000.00      1
 .664945270E+01 .226232110E-01-.806420670E-05 .954149200E-09 .000000000E+00    2
 .206794519E+05-.786429084E+01 .283048200E+00 .386777000E-01-.210739710E-04    3
 .427582900E-08 .000000000E+00 .225247800E+05 .254564400E+02                   4
RMP3                    C   4H   7O   2     G    300.00   4000.00 1376.00      1
 .154260382E+02 .169789201E-01-.593961909E-05 .936106835E-09-.548809672E-13    2
-.343012110E+05-.525677530E+02 .406577480E+01 .388324925E-01-.208048750E-04    3
 .506251249E-08-.421741752E-12-.297848227E+05 .102796868E+02                   4
NC4H9S                  C   4H   9          G    300.00   4000.00 1000.00      1
 .182440000E+01 .354350280E-01-.136901980E-04 .172985780E-08 .000000000E+00    2
 .521137543E+04 .190721830E+02 .882678800E+00 .419813690E-01-.239577090E-04    3
 .639274900E-08 .000000000E+00 .513670700E+04 .226104800E+02                   4
NC4H9P                  C   4H   9          G    300.00   4000.00 1000.00      1
 .285927140E+01 .339093470E-01-.129634890E-04 .162487360E-08 .000000000E+00    2
 .644131902E+04 .136765387E+02 .361027200E+00 .446560900E-01-.269622400E-04    3
 .737512580E-08 .000000000E+00 .679487900E+04 .252696800E+02                   4
IC4H9T                  C   4H   9          G    300.00   4000.00 1000.00      1
 .678309830E+01 .275756420E-01-.999251920E-05 .119923980E-08 .000000000E+00    2
 .130943964E+04-.110379681E+02-.668177200E+00 .478197410E-01-.281268890E-04    3
 .654078610E-08 .000000000E+00 .334806900E+04 .274761900E+02                   4
IC4H9P                  C   4H   9          G    300.00   4000.00 1000.00      1
 .672898190E+01 .277240280E-01-.100574610E-04 .120817530E-08 .000000000E+00    2
 .390175463E+04-.921990655E+01-.514098700E+00 .469939600E-01-.268680800E-04    3
 .599194290E-08 .000000000E+00 .591746700E+04 .283543100E+02                   4
CH3CH2CH2CHOH           C   4H   9O   1     G    300.00   4000.00 1389.00      1
 .146211284E+02 .192812832E-01-.662005863E-05 .103030580E-08-.598746774E-13    2
-.185860609E+05-.491894138E+02 .151231967E+01 .485940354E-01-.319829373E-04    3
 .112440534E-07-.168373464E-11-.138241933E+05 .218089522E+02                   4
CH3CHCH3CHOH            C   4H   9O   1     G    300.00   4000.00 1673.00      1
 .145354872E+02 .193544788E-01-.655352544E-05 .101052180E-08-.583473661E-13    2
-.195307842E+05-.500528678E+02 .524328525E+00 .528985884E-01-.379651080E-04    3
 .147054933E-07-.239054621E-11-.147012758E+05 .249822692E+02                   4
CH3CH2COHCH3            C   4H   9O   1     G    300.00   4000.00 1390.00      1
 .151619233E+02 .189741815E-01-.654734215E-05 .102237774E-08-.595503510E-13    2
-.208549516E+05-.532957109E+02 .108860217E+01 .524153990E-01-.380997951E-04    3
 .151074363E-07-.254404184E-11-.159195374E+05 .222613243E+02                   4
RTC4H8OH                C   4H   9O   1     G    300.00   4000.00 1395.00      1
 .146782533E+02 .193935063E-01-.660052048E-05 .102120044E-08-.590998119E-13    2
-.199408575E+05-.505292168E+02-.836665970E-01 .558040633E-01-.420184309E-04    3
 .171111519E-07-.290735214E-11-.149499995E+05 .281627857E+02                   4
RTC4H9O                 C   4H   9O   1     G    300.00   4000.00 1391.00      1
 .154820006E+02 .191120896E-01-.659337031E-05 .102954283E-08-.599712426E-13    2
-.189474281E+05-.587209701E+02-.652960434E+00 .575360662E-01-.423660204E-04    3
 .165461682E-07-.269335532E-11-.133634774E+05 .277645681E+02                   4
CH2CH2CHOHCH3           C   4H   9O   1     G    300.00   4000.00 1390.00      1
 .147487308E+02 .193476286E-01-.668165997E-05 .104395798E-08-.608330722E-13    2
-.178485397E+05-.492109234E+02 .467890397E+00 .521732276E-01-.362067190E-04    3
 .135025449E-07-.213961182E-11-.127480216E+05 .278224820E+02                   4
CH3CH2CHCH2OH           C   4H   9O   1     G    300.00   4000.00 2017.00      1
 .125195208E+02 .211308942E-01-.735078190E-05 .116027279E-08-.682567448E-13    2
-.159698333E+05-.352643597E+02 .927266773E+00 .453885784E-01-.244944451E-04    3
 .574420616E-08-.382704524E-12-.119074306E+05 .276532069E+02                   4
CH3CHCH2CH2OH           C   4H   9O   1     G    300.00   4000.00 2017.00      1
 .125195208E+02 .211308942E-01-.735078190E-05 .116027279E-08-.682567448E-13    2
-.159698333E+05-.352643597E+02 .927266773E+00 .453885784E-01-.244944451E-04    3
 .574420616E-08-.382704524E-12-.119074306E+05 .276532069E+02                   4
CH3CH2CHOHCH2           C   4H   9O   1     G    300.00   4000.00 1390.00      1
 .147487308E+02 .193476286E-01-.668165997E-05 .104395798E-08-.608330722E-13    2
-.178485397E+05-.492109234E+02 .467890397E+00 .521732276E-01-.362067190E-04    3
 .135025449E-07-.213961182E-11-.127480216E+05 .278224820E+02                   4
CH2CHCH2OHCH3           C   4H   9O   1     G    300.00   4000.00 1422.00      1
 .140854789E+02 .197806925E-01-.671026390E-05 .103599950E-08-.598718336E-13    2
-.165129917E+05-.457671006E+02-.566170728E-01 .523981203E-01-.356379876E-04    3
 .128198684E-07-.192264202E-11-.115334457E+05 .303769293E+02                   4
CH3CHCH2OCH3            C   4H   9O   1     G    300.00   4000.00 1422.00      1
 .148239632E+02 .195938055E-01-.674334212E-05 .105133556E-08-.611769464E-13    2
-.154937986E+05-.535942326E+02-.581327100E+00 .539666459E-01-.358338761E-04    3
 .122179671E-07-.171024843E-11-.995421675E+04 .297619860E+02                   4
CH3CCH2OHCH3            C   4H   9O   1     G    300.00   4000.00 1682.00      1
 .125605997E+02 .210637488E-01-.715019648E-05 .110439262E-08-.638428695E-13    2
-.183183621E+05-.368996627E+02 .329612707E+01 .347649647E-01-.102505618E-04    3
-.204641931E-08 .118879408E-11-.142607619E+05 .157499123E+02                   4
CH3CH2CHOCH3            C   4H   9O   1     G    300.00   4000.00 1382.00      1
 .157118766E+02 .189436692E-01-.663728010E-05 .104718616E-08-.614402720E-13    2
-.169625442E+05-.584079611E+02-.123566480E+00 .537328693E-01-.359804830E-04    3
 .125064763E-07-.182873667E-11-.111514942E+05 .275750096E+02                   4
CH3CH2CH2CH2O           C   4H   9O   1     G    300.00   4000.00 1383.00      1
 .150639724E+02 .192754979E-01-.670246160E-05 .105215438E-08-.615166356E-13    2
-.145981078E+05-.535775104E+02 .266423313E+00 .503656318E-01-.308368147E-04    3
 .928122753E-08-.110203449E-11-.905887861E+04 .272172881E+02                   4
CH3CHCHOHCH3            C   4H   9O   1     G    300.00   4000.00 1387.00      1
 .142049192E+02 .195897318E-01-.671801693E-05 .104483881E-08-.606940644E-13    2
-.190416934E+05-.463876157E+02 .933300006E+00 .472805232E-01-.278316313E-04    3
 .797039080E-08-.870532264E-12-.140666468E+05 .261224696E+02                   4
CH2CH2CH2CH2OH          C   4H   9O   1     G    300.00   4000.00 1388.00      1
 .142154423E+02 .196229836E-01-.673796562E-05 .104876785E-08-.609536943E-13    2
-.155756339E+05-.451352578E+02 .916505889E+00 .482692226E-01-.299841815E-04    3
 .956515610E-08-.126002465E-11-.106572242E+05 .272437766E+02                   4
NC4-QOOH                C   4H   9O   2     G    300.00   4000.00 1391.00      1
 .182943014E+02 .184250091E-01-.627217889E-05 .971379578E-09-.562825607E-13    2
-.128564704E+05-.650917535E+02 .986162058E+00 .585630676E-01-.416710545E-04    3
 .151223447E-07-.222454695E-11-.684048054E+04 .279289603E+02                   4
NC4H9-OO                C   4H   9O   2     G    300.00   4000.00 1392.00      1
 .164199470E+02 .207668293E-01-.714061871E-05 .111233445E-08-.646799300E-13    2
-.172909027E+05-.576444825E+02 .859225542E+00 .589774363E-01-.445935184E-04    3
 .184502497E-07-.321329944E-11-.119598721E+05 .254554544E+02                   4
IC4T-QOOH               C   4H   9O   2     G    300.00   4000.00 1397.00      1
 .188631296E+02 .183239932E-01-.631233086E-05 .984688082E-09-.573186521E-13    2
-.138981290E+05-.708829284E+02-.425033602E+00 .698121411E-01-.606175877E-04    3
 .274812344E-07-.501908797E-11-.779203954E+04 .305104370E+02                   4
IC4P-QOOH               C   4H   9O   2     G    300.00   4000.00 1396.00      1
 .181457399E+02 .188972595E-01-.650258715E-05 .101363925E-08-.589752496E-13    2
-.103249571E+05-.654833345E+02-.253900783E+00 .658110437E-01-.535280232E-04    3
 .228723790E-07-.398637599E-11-.429699727E+04 .319918975E+02                   4
IC4H9T-OO               C   4H   9O   2     G    300.00   4000.00 1392.00      1
 .167547908E+02 .205266172E-01-.706765238E-05 .110199004E-08-.641203511E-13    2
-.197490954E+05-.625129056E+02 .429458545E+00 .619305024E-01-.492178248E-04    3
 .213391061E-07-.385156685E-11-.142778206E+05 .242205126E+02                   4
IC4H9P-OO               C   4H   9O   2     G    300.00   4000.00 1391.00      1
 .160321835E+02 .211162441E-01-.726598082E-05 .113244436E-08-.658740064E-13    2
-.161760498E+05-.559920048E+02 .591660961E+00 .579744782E-01-.422019324E-04    3
 .167841571E-07-.283252682E-11-.107815683E+05 .268393730E+02                   4
RBU1OOX                 C   4H   9O   3     G    300.00   4000.00 1392.00      1
 .179101133E+02 .211247449E-01-.724787505E-05 .112742547E-08-.654930094E-13    2
-.371878276E+05-.612769774E+02 .289779336E+01 .560720331E-01-.390996379E-04    3
 .147174953E-07-.234862827E-11-.318812119E+05 .195265598E+02                   4
QBU1OOX                 C   4H   9O   3     G    300.00   4000.00 1386.00      1
 .129455763E+02 .795235476E-02-.280679691E-05 .445205248E-09-.262240810E-13    2
 .175946397E+05-.478819894E+02-.584674088E+01 .620875882E-01-.630010605E-04    3
 .306882361E-07-.575456234E-11 .230253176E+05 .492940922E+02                   4
IC4T-OOQOOH             C   4H   9O   4     G    300.00   4000.00 1391.00      1
 .225796674E+02 .201772761E-01-.702773819E-05 .110438266E-08-.646157968E-13    2
-.320684788E+05-.852469773E+02 .152317721E+01 .757827720E-01-.656981278E-04    3
 .300159936E-07-.556277284E-11-.252715176E+05 .257762885E+02                   4
IC4P-OOQOOH             C   4H   9O   4     G    300.00   4000.00 1390.00      1
 .218612263E+02 .207812365E-01-.723484570E-05 .113659545E-08-.664871920E-13    2
-.284979533E+05-.798472350E+02 .156900216E+01 .724191880E-01-.596183448E-04    3
 .260680737E-07-.468228506E-11-.217597632E+05 .278260039E+02                   4
NC4-OOQOOH              C   4H   9O   4     G    300.00   4000.00 1393.00      1
 .231119306E+02 .196469811E-01-.682730172E-05 .107124796E-08-.626109519E-13    2
-.320261199E+05-.872192509E+02 .109604492E+01 .794472856E-01-.714221316E-04    3
 .334124791E-07-.626730135E-11-.251118713E+05 .282288973E+02                   4
ZBU1OOX                 C   4H   9O   5     G    300.00   4000.00 1397.00      1
 .236719411E+02 .205751255E-01-.708127339E-05 .110392970E-08-.642301320E-13    2
-.515463449E+05-.860806755E+02 .475209184E+01 .678608013E-01-.534336966E-04    3
 .221852722E-07-.378003417E-11-.452511232E+05 .144907043E+02                   4
CYC5H5                  C   5H   5          G    300.00   4000.00 1000.00      1
 .421464919E+01 .271834728E-01-.133173209E-04 .308980119E-08-.277879873E-12    2
 .288952416E+05-.305999781E-01-.737844042E+01 .972391818E-01-.169579138E-03    3
 .151818667E-06-.512075479E-10 .305514662E+05 .512829539E+02                   4
C5H5O                   C   5H   5O   1     G    300.00   4000.00 1395.00      1
 .149072105E+02 .136369619E-01-.470762207E-05 .736028654E-09-.429314124E-13    2
 .143724130E+05-.569296345E+02-.414628450E+01 .623584874E-01-.528374678E-04    3
 .224628793E-07-.380136191E-11 .204992627E+05 .437921058E+02                   4
C5H7                    C   5H   7          G    300.00   4000.00 1000.00      1
 .671323690E+01 .274278890E-01-.994311090E-05 .119373240E-08 .000000000E+00    2
 .235116384E+05-.112735252E+02 .759315300E+00 .432678800E-01-.237613290E-04    3
 .512588110E-08 .000000000E+00 .251686000E+05 .196131100E+02                   4
RMCROTA                 C   5H   7O   2     G    300.00   4000.00 1000.00      1
 .151681730E+02 .178142000E-01-.496258460E-05 .688767770E-09-.386765100E-13    2
-.320532540E+05-.462913590E+02-.242828070E+00 .630479530E-01-.556979940E-04    3
 .265678430E-07-.501508770E-11-.278218120E+05 .329157640E+02                   4
NC5H9                   C   5H   9          G    300.00   4000.00 1383.00      1
 .140838604E+02 .208584950E-01-.722620456E-05 .113154433E-08-.660424465E-13    2
 .542225436E+04-.515371079E+02-.697079542E+00 .514354766E-01-.304500502E-04    3
 .880925852E-08-.994458078E-12 .110172568E+05 .293601364E+02                   4
NC5H9-5                 C   5H   9          G    300.00   4000.00 1383.00      1
 .140838604E+02 .208584950E-01-.722620456E-05 .113154433E-08-.660424465E-13    2
 .542225436E+04-.515371079E+02-.697079542E+00 .514354766E-01-.304500502E-04    3
 .880925852E-08-.994458078E-12 .110172568E+05 .293601364E+02                   4
NC5H9-4                 C   5H   9          G    300.00   4000.00 1383.00      1
 .140838604E+02 .208584950E-01-.722620456E-05 .113154433E-08-.660424465E-13    2
 .542225436E+04-.515371079E+02-.697079542E+00 .514354766E-01-.304500502E-04    3
 .880925852E-08-.994458078E-12 .110172568E+05 .293601364E+02                   4
NC5H9-3                 C   5H   9          G    300.00   4000.00 1383.00      1
 .140838604E+02 .208584950E-01-.722620456E-05 .113154433E-08-.660424465E-13    2
 .542225436E+04-.515371079E+02-.697079542E+00 .514354766E-01-.304500502E-04    3
 .880925852E-08-.994458078E-12 .110172568E+05 .293601364E+02                   4
C5EN-QOOH-43            C   5H   9O   2     G    300.00   4000.00 1392.00      1
 .203810644E+02 .199415880E-01-.695158032E-05 .109308002E-08-.639829228E-13    2
-.198146484E+02-.759778447E+02 .111814871E+01 .671698903E-01-.526574214E-04    3
 .218036776E-07-.373297383E-11 .652627032E+04 .268196384E+02                   4
C5EN-OO-4               C   5H   9O   2     G    300.00   4000.00 1392.00      1
 .186695690E+02 .216228347E-01-.748565666E-05 .117148772E-08-.683420517E-13    2
-.458976288E+04-.678082548E+02 .338814185E+00 .676913346E-01-.538434525E-04    3
 .231725654E-07-.414643363E-11 .158489053E+04 .297116190E+02                   4
C5EN-QOOH-34            C   5H   9O   2     G    300.00   4000.00 1392.00      1
 .203810644E+02 .199415880E-01-.695158032E-05 .109308002E-08-.639829228E-13    2
-.198146484E+02-.759778447E+02 .111814871E+01 .671698903E-01-.526574214E-04    3
 .218036776E-07-.373297383E-11 .652627032E+04 .268196384E+02                   4
C5EN-QOOH-35            C   5H   9O   2     G    300.00   4000.00 1392.00      1
 .203810644E+02 .199415880E-01-.695158032E-05 .109308002E-08-.639829228E-13    2
-.198146484E+02-.759778447E+02 .111814871E+01 .671698903E-01-.526574214E-04    3
 .218036776E-07-.373297383E-11 .652627032E+04 .268196384E+02                   4
C5EN-OO-3               C   5H   9O   2     G    300.00   4000.00 1392.00      1
 .186695690E+02 .216228347E-01-.748565666E-05 .117148772E-08-.683420517E-13    2
-.458976288E+04-.678082548E+02 .338814185E+00 .676913346E-01-.538434525E-04    3
 .231725654E-07-.414643363E-11 .158489053E+04 .297116190E+02                   4
C5EN-OO-5               C   5H   9O   2     G    300.00   4000.00 1392.00      1
 .186695690E+02 .216228347E-01-.748565666E-05 .117148772E-08-.683420517E-13    2
-.458976288E+04-.678082548E+02 .338814185E+00 .676913346E-01-.538434525E-04    3
 .231725654E-07-.414643363E-11 .158489053E+04 .297116190E+02                   4
RMBX                    C   5H   9O   2     G    300.00   4000.00 1382.00      1
 .193382201E+02 .209401493E-01-.732209753E-05 .115371679E-08-.676297088E-13    2
-.412852468E+05-.755834444E+02 .231680806E+01 .569247905E-01-.356059275E-04    3
 .110212330E-07-.136558032E-11-.349304634E+05 .172843303E+02                   4
C5EN-QOOH-53            C   5H   9O   2     G    300.00   4000.00 1392.00      1
 .203810644E+02 .199415880E-01-.695158032E-05 .109308002E-08-.639829228E-13    2
-.198146484E+02-.759778447E+02 .111814871E+01 .671698903E-01-.526574214E-04    3
 .218036776E-07-.373297383E-11 .652627032E+04 .268196384E+02                   4
C5EN-QOOH-45            C   5H   9O   2     G    300.00   4000.00 1392.00      1
 .203810644E+02 .199415880E-01-.695158032E-05 .109308002E-08-.639829228E-13    2
-.198146484E+02-.759778447E+02 .111814871E+01 .671698903E-01-.526574214E-04    3
 .218036776E-07-.373297383E-11 .652627032E+04 .268196384E+02                   4
C5EN-QOOH-54            C   5H   9O   2     G    300.00   4000.00 1392.00      1
 .203810644E+02 .199415880E-01-.695158032E-05 .109308002E-08-.639829228E-13    2
-.198146484E+02-.759778447E+02 .111814871E+01 .671698903E-01-.526574214E-04    3
 .218036776E-07-.373297383E-11 .652627032E+04 .268196384E+02                   4
C5EN-OOQOOH-43          C   5H   9O   4     G    300.00   4000.00 1000.00      1
 .251889054E+02 .206642290E-01-.723193822E-05 .114017997E-08-.668636462E-13    2
-.189404232E+05-.976775550E+02 .705279661E+00 .861579519E-01-.769448689E-04    3
 .356373390E-07-.663192053E-11-.111524362E+05 .310665731E+02                   4
C5EN-OOQOOH-34          C   5H   9O   4     G    300.00   4000.00 1000.00      1
 .251889054E+02 .206642290E-01-.723193822E-05 .114017997E-08-.668636462E-13    2
-.189404232E+05-.976775550E+02 .705279661E+00 .861579519E-01-.769448689E-04    3
 .356373390E-07-.663192053E-11-.111524362E+05 .310665731E+02                   4
QMBOOX                  C   5H   9O   4     G    300.00   4000.00 1000.00      1
 .211938570E+02 .222144000E-01-.631327380E-05 .888168590E-09-.502931100E-13    2
-.572489530E+05-.734085620E+02 .256566330E+01 .606897660E-01-.678613150E-05    3
-.390168040E-07 .205529000E-10-.518452190E+05 .251823650E+02                   4
RMBOOX                  C   5H   9O   4     G    300.00   4000.00 1000.00      1
 .211938570E+02 .222144000E-01-.631327380E-05 .888168590E-09-.502931100E-13    2
-.572489530E+05-.734085620E+02 .256566330E+01 .606897660E-01-.678613150E-05    3
-.390168040E-07 .205529000E-10-.518452190E+05 .251823650E+02                   4
C5EN-OOQOOH-53          C   5H   9O   4     G    300.00   4000.00 1000.00      1
 .251889054E+02 .206642290E-01-.723193822E-05 .114017997E-08-.668636462E-13    2
-.189404232E+05-.976775550E+02 .705279661E+00 .861579519E-01-.769448689E-04    3
 .356373390E-07-.663192053E-11-.111524362E+05 .310665731E+02                   4
C5EN-OOQOOH-45          C   5H   9O   4     G    300.00   4000.00 1000.00      1
 .251889054E+02 .206642290E-01-.723193822E-05 .114017997E-08-.668636462E-13    2
-.189404232E+05-.976775550E+02 .705279661E+00 .861579519E-01-.769448689E-04    3
 .356373390E-07-.663192053E-11-.111524362E+05 .310665731E+02                   4
C5EN-OOQOOH-35          C   5H   9O   4     G    300.00   4000.00 1000.00      1
 .251889054E+02 .206642290E-01-.723193822E-05 .114017997E-08-.668636462E-13    2
-.189404232E+05-.976775550E+02 .705279661E+00 .861579519E-01-.769448689E-04    3
 .356373390E-07-.663192053E-11-.111524362E+05 .310665731E+02                   4
C5EN-OOQOOH-54          C   5H   9O   4     G    300.00   4000.00 1000.00      1
 .251889054E+02 .206642290E-01-.723193822E-05 .114017997E-08-.668636462E-13    2
-.189404232E+05-.976775550E+02 .705279661E+00 .861579519E-01-.769448689E-04    3
 .356373390E-07-.663192053E-11-.111524362E+05 .310665731E+02                   4
ZMBOOX                  C   5H   9O   6     G    300.00   4000.00 1000.00      1
 .261471200E+02 .215283560E-01-.581135510E-05 .785452200E-09-.431572980E-13    2
-.689643590E+05-.913329620E+02 .443715430E+01 .699071290E-01-.165602940E-04    3
-.356586160E-07 .205531550E-10-.628690510E+05 .226288070E+02                   4
NC5H11                  C   5H  11          G    300.00   4000.00 1384.00      1
 .131340658E+02 .260923466E-01-.897731137E-05 .139920325E-08-.813970860E-13    2
-.427735231E+04-.434455998E+02-.304386354E+01 .581995422E-01-.316090839E-04    3
 .790004927E-08-.665198232E-12 .199185425E+04 .455946950E+02                   4
NEOC5H11                C   5H  11          G    300.00   4000.00 1396.00      1
 .166235914E+02 .227037884E-01-.771624835E-05 .119289853E-08-.690060600E-13    2
-.396429146E+04-.644693953E+02-.158140132E+01 .657175067E-01-.468120314E-04    3
 .174732793E-07-.268709925E-11 .230933742E+04 .331296742E+02                   4
C5H10-OH                C   5H  11O   1     G    300.00   4000.00 1392.00      1
 .199150940E+02 .250390538E-01-.861981469E-05 .134386616E-08-.781893344E-13    2
-.238472344E+05-.769667628E+02 .235935841E+00 .739755736E-01-.572379508E-04    3
 .241234657E-07-.425357119E-11-.171710700E+05 .279024996E+02                   4
RMTBE                   C   5H  11O   1     G    300.00   4000.00 1386.00      1
 .191923401E+02 .226496418E-01-.770522799E-05 .119249279E-08-.690514122E-13    2
-.223486482E+05-.717004889E+02-.284403552E+00 .706092470E-01-.543641242E-04    3
 .224557925E-07-.385680161E-11-.157511970E+05 .321647207E+02                   4
NEOC5H11-OO             C   5H  11O   2     G    300.00   4000.00 1396.00      1
 .202154849E+02 .245786365E-01-.841704919E-05 .130775217E-08-.759095109E-13    2
-.224777899E+05-.796085899E+02 .730403748E+00 .705036948E-01-.502866599E-04    3
 .189083885E-07-.294948183E-11-.157211898E+05 .249439750E+02                   4
NC5-QOOH                C   5H  11O   2     G    300.00   4000.00 1396.00      1
 .220245928E+02 .228314385E-01-.786198359E-05 .122609365E-08-.713571493E-13    2
-.179960313E+05-.864387261E+02-.607426660E+00 .818016374E-01-.685494236E-04    3
 .302071532E-07-.540750321E-11-.106868081E+05 .330450153E+02                   4
NC5H12OO                C   5H  11O   2     G    300.00   4000.00 1392.00      1
 .199150940E+02 .250390538E-01-.861981469E-05 .134386616E-08-.781893344E-13    2
-.238472344E+05-.769667628E+02 .235935841E+00 .739755736E-01-.572379508E-04    3
 .241234657E-07-.425357119E-11-.171710700E+05 .279024996E+02                   4
NEOC5-QOOH              C   5H  11O   2     G    300.00   4000.00 1396.00      1
 .218550366E+02 .228989820E-01-.786956915E-05 .122572909E-08-.712760383E-13    2
-.164801773E+05-.857429310E+02 .115441893E+01 .724266160E-01-.535668095E-04    3
 .205704339E-07-.323425526E-11-.941504872E+04 .250054329E+02                   4
MTBE-OO                 C   5H  11O   3     G    300.00   4000.00 1386.00      1
 .219476262E+02 .253064866E-01-.877948807E-05 .137597948E-08-.803553517E-13    2
-.383949561E+05-.811182382E+02 .226233362E+01 .712292692E-01-.511734982E-04    3
 .199100134E-07-.329751069E-11-.314029562E+05 .248780910E+02                   4
MTBE-QOOH               C   5H  11O   3     G    300.00   4000.00 1401.00      1
 .214971173E+02 .259064341E-01-.848605930E-05 .127921441E-08-.726936886E-13    2
-.312441531E+05-.765479844E+02 .134883146E+01 .795292274E-01-.643595941E-04    3
 .280404405E-07-.497823206E-11-.249060790E+05 .293286141E+02                   4
C5H10-OHOO              C   5H  11O   3     G    300.00   4000.00 1392.00      1
 .199150940E+02 .250390538E-01-.861981469E-05 .134386616E-08-.781893344E-13    2
-.238472344E+05-.769667628E+02 .235935841E+00 .739755736E-01-.572379508E-04    3
 .241234657E-07-.425357119E-11-.171710700E+05 .279024996E+02                   4
NC5-OOQOOH              C   5H  11O   4     G    300.00   4000.00 1391.00      1
 .257270270E+02 .247172056E-01-.859292907E-05 .134865114E-08-.788382618E-13    2
-.361631686E+05-.100728579E+03 .135798731E+01 .877212925E-01-.735867140E-04    3
 .327395450E-07-.595540146E-11-.281695250E+05 .282261555E+02                   4
NEOC5-OOQOOH            C   5H  11O   4     G    300.00   4000.00 1392.00      1
 .248490803E+02 .252599638E-01-.873651764E-05 .136662251E-08-.797082603E-13    2
-.350133010E+05-.961825156E+02 .265748524E+01 .758789336E-01-.526594216E-04    3
 .186692316E-07-.269820831E-11-.271776626E+05 .234450387E+02                   4
MTBE-OOQOOH             C   5H  11O   5     G    300.00   4000.00 1391.00      1
 .264681284E+02 .261757287E-01-.899393547E-05 .140058534E-08-.814301239E-13    2
-.504985383E+05-.992053288E+02 .454595241E+01 .801871705E-01-.616423289E-04    3
 .254521416E-07-.437448229E-11-.430642384E+05 .177072264E+02                   4
C6H3                    C   6H   3          G    300.00   4000.00 1000.00      1
 .120132339E+02 .114461128E-01-.408884040E-05 .657753914E-09-.392832116E-13    2
 .825892145E+05-.335118700E+02 .150089155E+01 .545901804E-01-.788221454E-04    3
 .627969099E-07-.200768594E-10 .849133510E+05 .176237455E+02                   4
LC6H5                   C   6H   5          G    300.00   4000.00 1000.00      1
 .134117680E+02 .147202210E-01-.508177050E-05 .798863540E-09-.469508440E-13    2
 .585037160E+05-.416520320E+02 .779297070E+00 .543721260E-01-.478738140E-04    3
 .161871640E-07 .337357440E-12 .616503120E+05 .221285920E+02                   4
C6H5                    C   6H   5          G    300.00   4000.00 1000.00      1
 .157758892E+02 .965110900E-02-.942941600E-06-.546911100E-09 .102652200E-12    2
 .330269797E+05-.617628096E+02 .114355700E+00 .362732400E-01 .115828600E-05    3
-.219696400E-07 .846355600E-11 .383605400E+05 .238011700E+02                   4
C6H5O                   C   6H   5O   1     G    300.00   4000.00 1000.00      1
 .137221720E+02 .174688771E-01-.635504520E-05 .103492308E-08-.623410504E-13    2
 .287274751E+03-.488181680E+02-.466204455E+00 .413443975E-01 .132412991E-04    3
-.572872769E-07 .289763707E-10 .477858391E+04 .276990274E+02                   4
DMF-3YL                 C   6H   7O   1     G    300.00   4000.00 1000.00      1
 .118002735E+02 .257930235E-01-.101089409E-04 .181299326E-08-.122176870E-12    2
 .130508362E+05-.352008048E+02 .197118616E+01 .384836786E-01 .786460722E-05    3
-.354301012E-07 .162325679E-10 .165648455E+05 .193223377E+02                   4
CYC6H9                  C   6H   9          G    300.00   4000.00 1381.00      1
 .166730638E+02 .227088190E-01-.801509353E-05 .127088484E-08-.748275111E-13    2
 .698387216E+04-.723601536E+02-.631908086E+01 .726795534E-01-.484456826E-04    3
 .157628084E-07-.202092558E-11 .153574632E+05 .524769640E+02                   4
RALDEST                 C   6H   9O   3     G    300.00   4000.00 1373.00      1
 .215153215E+02 .236419666E-01-.830694270E-05 .131026314E-08-.767602984E-13    2
-.530993462E+05-.770487448E+02 .687062608E+01 .492844450E-01-.217786396E-04    3
 .243527207E-08 .464021620E-12-.470662293E+05 .479532953E+01                   4
CYC6H11                 C   6H  11          G    300.00   4000.00 1674.00      1
 .146799252E+02 .309324453E-01-.112934485E-04 .183887582E-08-.110464203E-12    2
-.197594614E+03-.590168221E+02-.757310296E+01 .766896480E-01-.424441426E-04    3
 .941423236E-08-.439999709E-12 .764576045E+04 .620172120E+02                   4
CYC6-QOOH-2             C   6H  11O   2     G    300.00   4000.00 1375.00      1
 .243899542E+02 .262326944E-01-.930434909E-05 .148019558E-08-.873538395E-13    2
-.163135893E+05-.107549099E+03-.378907832E+01 .841562901E-01-.510965662E-04    3
 .133666762E-07-.102528616E-11-.580881865E+04 .464783226E+02                   4
CYC6-QOOH-3             C   6H  11O   2     G    300.00   4000.00 1374.00      1
 .241250295E+02 .262273012E-01-.925328534E-05 .146724451E-08-.864028312E-13    2
-.163808524E+05-.106267870E+03-.596804450E+01 .893075551E-01-.558813589E-04    3
 .152003723E-07-.125762311E-11-.534935832E+04 .576800888E+02                   4
CYC6-OO                 C   6H  11O   2     G    300.00   4000.00 1380.00      1
 .225527144E+02 .280656231E-01-.990087442E-05 .156942170E-08-.923867180E-13    2
-.209455781E+05-.994788807E+02-.594021024E+01 .887171975E-01-.569424328E-04    3
 .171601250E-07-.191055830E-11-.104841379E+05 .556048484E+02                   4
CYC6-QOOH-4             C   6H  11O   2     G    300.00   4000.00 1374.00      1
 .241250295E+02 .262273012E-01-.925328534E-05 .146724451E-08-.864028312E-13    2
-.163808524E+05-.106267870E+03-.596804450E+01 .893075551E-01-.558813589E-04    3
 .152003723E-07-.125762311E-11-.534935832E+04 .576800888E+02                   4
CYC6-OOQOOH-4           C   6H  11O   4     G    300.00   4000.00 1383.00      1
 .291238921E+02 .270060308E-01-.959994599E-05 .152947435E-08-.903544360E-13    2
-.353659440E+05-.128893429E+03-.534585270E+01 .106448443E+00-.790742157E-04    3
 .290275771E-07-.426034434E-11-.233396667E+05 .565320100E+02                   4
CYC6-OOQOOH-2           C   6H  11O   4     G    300.00   4000.00 1383.00      1
 .291238921E+02 .270060308E-01-.959994599E-05 .152947435E-08-.903544360E-13    2
-.353659440E+05-.128198915E+03-.534585270E+01 .106448443E+00-.790742157E-04    3
 .290275771E-07-.426034434E-11-.233396667E+05 .572265244E+02                   4
CYC6-OOQOOH-3           C   6H  11O   4     G    300.00   4000.00 1383.00      1
 .291238921E+02 .270060308E-01-.959994599E-05 .152947435E-08-.903544360E-13    2
-.353659440E+05-.128198915E+03-.534585270E+01 .106448443E+00-.790742157E-04    3
 .290275771E-07-.426034434E-11-.233396667E+05 .572265244E+02                   4
RDIPE                   C   6H  13O   1     G    300.00   4000.00 1389.00      1
 .195346832E+02 .300586517E-01-.103564671E-04 .161544621E-08-.940217507E-13    2
-.289625035E+05-.700231442E+02-.545711430E-01 .748436725E-01-.509801332E-04    3
 .191769721E-07-.313046382E-11-.218696353E+05 .358513387E+02                   4
C7H7                    C   7H   7          G    300.00   4000.00 1000.00      1
 .126890424E+02 .248754040E-01-.820402330E-05 .901804910E-09 .000000000E+00    2
 .179417186E+05-.454264236E+02-.296228400E+01 .659171040E-01-.433334430E-04    3
 .106408510E-07 .000000000E+00 .223472400E+05 .359657700E+02                   4
C6H4CH3                 C   7H   7          G    300.00   4000.00 1000.00      1
 .989521100E+01 .281997140E-01-.985390310E-05 .114532240E-08 .000000000E+00    2
 .307512908E+05-.257557742E+02-.298827000E+01 .621039310E-01-.390118950E-04    3
 .928257830E-08 .000000000E+00 .343676800E+05 .412025200E+02                   4
RCRESOLC                C   7H   7O   1     G    300.00   4000.00 1000.00      1
 .689970000E+01 .376640500E-01-.142499000E-04 .245139600E-08-.159215300E-12    2
-.104378100E+04-.796692700E+01-.415304900E+01 .776998800E-01-.583028700E-04    3
 .178677900E-07-.536299700E-12 .896696700E+03 .453288900E+02                   4
RCRESOLO                C   7H   7O   1     G    300.00   4000.00 1000.00      1
 .632623400E+01 .370920700E-01-.137369600E-04 .232847100E-08-.149701800E-12    2
-.156635900E+04-.468621100E+01-.403964400E+01 .739909500E-01-.515945300E-04    3
 .120372800E-07 .143210200E-11 .225707600E+03 .453169300E+02                   4
NC7H13                  C   7H  13          G    300.00   4000.00 1383.00      1
 .140838604E+02 .208584950E-01-.722620456E-05 .113154433E-08-.660424465E-13    2
 .542225436E+04-.515371079E+02-.697079542E+00 .514354766E-01-.304500502E-04    3
 .880925852E-08-.994458078E-12 .110172568E+05 .293601364E+02                   4
RMCYC6                  C   7H  13          G    300.00   4000.00 2030.00      1
 .173202469E+02 .361144629E-01-.130438584E-04 .210911191E-08-.126098895E-12    2
-.514813032E+04-.717714814E+02-.853970231E+01 .919151844E-01-.546389770E-04    3
 .144889205E-07-.127842414E-11 .374687760E+04 .679730355E+02                   4
RMCYC6-OO               C   7H  13O   2     G    300.00   4000.00 1386.00      1
 .252650839E+02 .325458915E-01-.113494502E-04 .178540172E-08-.104551384E-12    2
-.262255150E+05-.112686720E+03-.606776148E+01 .998265984E-01-.637962761E-04    3
 .191011484E-07-.207496071E-11-.148337709E+05 .575547331E+02                   4
MCYC6T-QOOH             C   7H  13O   2     G    300.00   4000.00 2055.00      1
 .234331685E+02 .347621964E-01-.124048044E-04 .199225952E-08-.118633947E-12    2
-.195868561E+05-.990888361E+02-.694095755E+01 .104651350E+00-.698281467E-04    3
 .219897276E-07-.260222584E-11-.958151058E+04 .634587763E+02                   4
NC7H13O2                C   7H  13O   2     G    300.00   4000.00 1383.00      1
 .140838604E+02 .208584950E-01-.722620456E-05 .113154433E-08-.660424465E-13    2
 .542225436E+04-.515371079E+02-.697079542E+00 .514354766E-01-.304500502E-04    3
 .880925852E-08-.994458078E-12 .110172568E+05 .293601364E+02                   4
MCYC6-QOOH              C   7H  13O   2     G    300.00   4000.00 2055.00      1
 .234331685E+02 .347621964E-01-.124048044E-04 .199225952E-08-.118633947E-12    2
-.195868561E+05-.990888361E+02-.694095755E+01 .104651350E+00-.698281467E-04    3
 .219897276E-07-.260222584E-11-.958151058E+04 .634587763E+02                   4
MCYC6-OOQOOH            C   7H  13O   4     G    300.00   4000.00 1394.00      1
 .305321225E+02 .326136355E-01-.113442944E-04 .178165385E-08-.104214977E-12    2
-.403458401E+05-.135302325E+03-.434829022E+01 .112403701E+00-.796910207E-04    3
 .277878216E-07-.380650779E-11-.281870009E+05 .524217373E+02                   4
MCYC6T-OOQOOH           C   7H  13O   4     G    300.00   4000.00 1394.00      1
 .305321225E+02 .326136355E-01-.113442944E-04 .178165385E-08-.104214977E-12    2
-.403458401E+05-.135302325E+03-.434829022E+01 .112403701E+00-.796910207E-04    3
 .277878216E-07-.380650779E-11-.281870009E+05 .524217373E+02                   4
NC7H15                  C   7H  15          G    300.00   4000.00 1382.00      1
 .216371448E+02 .323324804E-01-.109273807E-04 .168357060E-08-.971774091E-13    2
-.105877217E+05-.852228493E+02-.379155767E-01 .756726570E-01-.407473634E-04    3
 .932678943E-08-.492360745E-12-.235605303E+04 .337321506E+02                   4
NC7H15-OO               C   7H  15O   2     G    300.00   4000.00 1393.00      1
 .272928290E+02 .327034748E-01-.112483701E-04 .175282538E-08-.101955579E-12    2
-.235449480E+05-.109307876E+03 .137396160E+01 .925294066E-01-.644403647E-04    3
 .235223293E-07-.356678305E-11-.144154775E+05 .302419431E+02                   4
NC7-QOOH                C   7H  15O   2     G    300.00   4000.00 1000.00      1
 .449365222E+02 .384325070E-02-.181753210E-06-.116055420E-10 .168632530E-14    2
-.301866739E+05-.207157897E+03 .169959950E+01 .943723540E-01-.755904260E-04    3
 .401131540E-07-.120065810E-10-.147076150E+05 .283145640E+02                   4
NC7-OOQOOH              C   7H  15O   4     G    300.00   4000.00 1395.00      1
 .269436049E+02 .351661203E-01-.120111248E-04 .186268617E-08-.107974911E-12    2
-.478858130E+05-.104588181E+03 .234060326E+01 .923428863E-01-.637138459E-04    3
 .236026902E-07-.368902757E-11-.392112217E+05 .278171493E+02                   4
C6H4C2H                 C   8H   5          G    300.00   4000.00 1000.00      1
 .286860656E+02-.138698600E-01 .227211900E-04-.998822700E-08 .140859000E-11    2
 .560473490E+05-.127502636E+03-.293242200E+01 .660436800E-01-.395005000E-04    3
-.318303810E-08 .853003870E-11 .653240430E+05 .380586850E+02                   4
C6H5C2H2                C   8H   7          G    300.00   4000.00 1394.00      1
 .187667289E+02 .200619262E-01-.690883699E-05 .107799789E-08-.627759176E-13    2
 .376789029E+05-.760287256E+02-.272251268E+01 .709701368E-01-.527526320E-04    3
 .197369835E-07-.295890798E-11 .450007235E+05 .390143531E+02                   4
C8H9                    C   8H   9          G    300.00   4000.00 1000.00      1
 .179749910E+02 .239625180E-01-.715492520E-05 .103757720E-08-.596944840E-13    2
 .194242850E+05-.693345570E+02-.526520200E+01 .889877600E-01-.754492360E-04    3
 .341497320E-07-.666954430E-11 .259605610E+05 .509400020E+02                   4
RXYLENE                 C   8H   9          G    300.00   4000.00 1000.00      1
 .808697123E+01 .442230490E-01-.196920930E-04 .391313300E-08-.286780230E-12    2
 .152828351E+05-.180507988E+02-.244083000E+01 .750206000E-01-.520941000E-04    3
 .184357000E-07-.267709000E-11 .180599500E+05 .358328500E+02                   4
RUME7                   C   8H  13O   2     G    300.00   4000.00 1376.00      1
 .270534591E+02 .305004468E-01-.106520501E-04 .167796515E-08-.983020287E-13    2
-.363346010E+05-.107800076E+03 .366021323E+01 .765652941E-01-.421034444E-04    3
 .990005395E-08-.618141131E-12-.272971814E+05 .209764369E+02                   4
RME7                    C   8H  15O   2     G    300.00   4000.00 1382.00      1
 .283088733E+02 .346001847E-01-.117889297E-04 .182346779E-08-.105527368E-12    2
-.507031223E+05-.115791454E+03 .312712425E+01 .886538094E-01-.550709022E-04    3
 .172495936E-07-.218153163E-11-.414147165E+05 .212562509E+02                   4
IC8H17                  C   8H  17          G    300.00   4000.00 1000.00      1
 .210071027E+02 .400670210E-01-.122220840E-04 .179139180E-08-.103364050E-12    2
-.156827594E+05-.841376688E+02-.142527150E+01 .952433870E-01-.515412500E-04    3
 .269038680E-08 .557281520E-11-.909216410E+04 .335841900E+02                   4
IC8H17-OO               C   8H  17O   2     G    300.00   4000.00 1397.00      1
 .307492955E+02 .368544999E-01-.126522533E-04 .196915974E-08-.114442369E-12    2
-.380116818E+05-.129042218E+03-.126574300E+01 .113828908E+00-.844050615E-04    3
 .328104935E-07-.525271208E-11-.270886887E+05 .421608430E+02                   4
IC8T-QOOH               C   8H  17O   2     G    300.00   4000.00 1400.00      1
 .323288504E+02 .354286616E-01-.121434812E-04 .188811322E-08-.109661472E-12    2
-.319868602E+05-.136609837E+03-.150530420E+01 .118500203E+00-.910186246E-04    3
 .362481173E-07-.587667874E-11-.206807572E+05 .436006519E+02                   4
IC8-QOOH                C   8H  17O   2     G    300.00   4000.00 1400.00      1
 .323288504E+02 .354286616E-01-.121434812E-04 .188811322E-08-.109661472E-12    2
-.319868602E+05-.136609837E+03-.150530420E+01 .118500203E+00-.910186246E-04    3
 .362481173E-07-.587667874E-11-.206807572E+05 .436006519E+02                   4
IC8-OOQOOH              C   8H  17O   4     G    300.00   4000.00 1398.00      1
 .362956073E+02 .372755603E-01-.128091685E-04 .199516372E-08-.116026947E-12    2
-.507708950E+05-.153592254E+03 .134208862E+01 .119507370E+00-.864939904E-04    3
 .319097725E-07-.475802942E-11-.387629197E+05 .338018650E+02                   4
INDENYL                 C   9H   7          G    300.00   4000.00 1389.00      1
 .210619876E+02 .219045968E-01-.772700080E-05 .122481766E-08-.721012249E-13    2
 .270100509E+05-.947705468E+02-.627808779E+01 .881610767E-01-.698280991E-04    3
 .280009421E-07-.454051640E-11 .362473103E+05 .511874555E+02                   4
RC9H11                  C   9H  11          G    300.00   4000.00 1385.00      1
 .227307929E+02 .291439937E-01-.101635526E-04 .159859987E-08-.935933623E-13    2
 .481056390E+04-.975266902E+02-.180604559E+01 .826070356E-01-.539943357E-04    3
 .177716542E-07-.237645289E-11 .137819561E+05 .357292291E+02                   4
C10H7                   C  10H   7          G    300.00   4000.00 1000.00      1
 .146529084E+02 .356159360E-01-.121796480E-04 .138747960E-08 .000000000E+00    2
 .405898415E+05-.575649187E+02-.631700500E+01 .913910790E-01-.608201990E-04    3
 .152228010E-07 .000000000E+00 .464268700E+05 .512234700E+02                   4
C10H7O                  C  10H   7O   1     G    300.00   4000.00 1387.00      1
 .252263199E+02 .234793777E-01-.827533154E-05 .131107385E-08-.771548491E-13    2
 .188945294E+04-.112699321E+03-.234081413E+01 .850055448E-01-.590412510E-04    3
 .195981954E-07-.248272174E-11 .116463286E+05 .362009562E+02                   4
RTETRALIN               C  10H  11          G    300.00   4000.00 1393.00      1
 .274897602E+02 .290231662E-01-.101643070E-04 .160474752E-08-.942455736E-13    2
 .498834588E+04-.134140516E+03-.103201226E+02 .112759920E+00-.777366610E-04    3
 .248527119E-07-.289510552E-11 .183518811E+05 .701782401E+02                   4
RTETRAOO                C  10H  11O   2     G    300.00   4000.00 1393.00      1
 .325696052E+02 .270322587E-01-.103226960E-04 .172977036E-08-.105947326E-12    2
-.797598133E+04-.153101057E+03-.133437809E+02 .139730780E+00-.110918062E-03    3
 .406822937E-07-.565600132E-11 .639529388E+04 .899902305E+02                   4
RDECALIN                C  10H  17          G    300.00   4000.00 1393.00      1
 .266885367E+02 .438181872E-01-.149997894E-04 .233096426E-08-.135354849E-12    2
-.142864228E+05-.128706101E+03-.137726588E+02 .134621624E+00-.905467076E-04    3
 .298633466E-07-.381482514E-11-.121358784E+02 .896659972E+02                   4
RODECA                  C  10H  17          G    300.00   4000.00 1393.00      1
 .266885367E+02 .438181872E-01-.149997894E-04 .233096426E-08-.135354849E-12    2
-.142864228E+05-.128706101E+03-.137726588E+02 .134621624E+00-.905467076E-04    3
 .298633466E-07-.381482514E-11-.121358784E+02 .896659972E+02                   4
RDECOO                  C  10H  17O   2     G    300.00   4000.00 1379.00      1
 .223721095E+02 .276799389E-01-.974217376E-05 .154194767E-08-.906767646E-13    2
-.211451384E+05-.984373555E+02-.491663898E+01 .836156703E-01-.498338842E-04    3
 .127483629E-07-.918573704E-12-.109593466E+05 .507734668E+02                   4
QDECOOH                 C  10H  17O   2     G    300.00   4000.00 1379.00      1
 .223721095E+02 .276799389E-01-.974217376E-05 .154194767E-08-.906767646E-13    2
-.211451384E+05-.984373555E+02-.491663898E+01 .836156703E-01-.498338842E-04    3
 .127483629E-07-.918573704E-12-.109593466E+05 .507734668E+02                   4
ZDECA                   C  10H  17O   4     G    300.00   4000.00 1379.00      1
 .223721095E+02 .276799389E-01-.974217376E-05 .154194767E-08-.906767646E-13    2
-.211451384E+05-.984373555E+02-.491663898E+01 .836156703E-01-.498338842E-04    3
 .127483629E-07-.918573704E-12-.109593466E+05 .507734668E+02                   4
NC10H19                 C  10H  19          G    300.00   4000.00 1383.00      1
 .140838604E+02 .208584950E-01-.722620456E-05 .113154433E-08-.660424465E-13    2
 .542225436E+04-.515371079E+02-.697079542E+00 .514354766E-01-.304500502E-04    3
 .880925852E-08-.994458078E-12 .110172568E+05 .293601364E+02                   4
NC10H21                 C  10H  21          G    300.00   4000.00 1385.00      1
 .314447580E+02 .452778532E-01-.153145696E-04 .236072411E-08-.136311835E-12    2
-.229702700E+05-.131435127E+03-.930536886E+00 .113137924E+00-.664034118E-04    3
 .183220872E-07-.177128003E-11-.109890165E+05 .451328034E+02                   4
NC10H21-OO              C  10H  21O   2     G    300.00   4000.00 1392.00      1
 .347424373E+02 .481682266E-01-.165183738E-04 .256870455E-08-.149189141E-12    2
-.416206773E+05-.145293449E+03 .109633829E+01 .123998092E+00-.822926235E-04    3
 .288935474E-07-.426829326E-11-.295195291E+05 .366210584E+02                   4
NC10-QOOH               C  10H  21O   2     G    300.00   4000.00 1392.00      1
 .364873664E+02 .456938220E-01-.154604572E-04 .238346695E-08-.137626430E-12    2
-.370093465E+05-.152798812E+03 .883511244E+00 .125360621E+00-.820308363E-04    3
 .270294818E-07-.354081617E-11-.243570772E+05 .395546233E+02                   4
NC10-OOQOOH             C  10H  21O   4     G    300.00   4000.00 1393.00      1
 .419701067E+02 .470326141E-01-.162065055E-04 .252885796E-08-.147242779E-12    2
-.568721943E+05-.179987435E+03 .270340236E+01 .134161981E+00-.884509572E-04    3
 .291143638E-07-.380678318E-11-.428023111E+05 .324857210E+02                   4
C10H6CH3                C  11H   9          G    300.00   4000.00 1387.00      1
 .241866524E+02 .287085863E-01-.100040198E-04 .157283341E-08-.920615442E-13    2
 .317595121E+05-.107209439E+03-.148986180E+01 .837301572E-01-.531437515E-04    3
 .161159556E-07-.183550466E-11 .411521411E+05 .324161445E+02                   4
C10H7CH2                C  11H   9          G    300.00   4000.00 1389.00      1
 .266596927E+02 .269903845E-01-.949827903E-05 .150313533E-08-.883831941E-13    2
 .210179470E+05-.122975754E+03-.551514480E+01 .106245066E+00-.857510752E-04    3
 .355122444E-07-.598055713E-11 .318146452E+05 .484291679E+02                   4
CH3C10H6O               C  11H   9O   1     G    300.00   4000.00 1386.00      1
 .281108749E+02 .281427040E-01-.986090177E-05 .155620703E-08-.913337710E-13    2
-.350666986E+04-.125748079E+03-.108570461E+01 .905308669E-01-.577474885E-04    3
 .167977934E-07-.168045736E-11 .709977655E+04 .329292729E+02                   4
RUME10                  C  11H  19O   2     G    300.00   4000.00 1400.00      1
 .333201898E+02 .479399831E-01-.157699228E-04 .238393079E-08-.135735725E-12    2
-.400970534E+05-.137405141E+03 .142231026E+01 .127120401E+00-.922642215E-04    3
 .364453822E-07-.599028369E-11-.294852312E+05 .322500169E+02                   4
RMDX                    C  11H  21O   2     G    300.00   4000.00 1376.00      1
 .385051195E+02 .464902832E-01-.162008540E-04 .254969816E-08-.149299808E-12    2
-.649901621E+05-.166525707E+03 .345128941E+01 .114960511E+00-.621890037E-04    3
 .140937438E-07-.752795690E-12-.513892174E+05 .266431624E+02                   4
RMDOOX                  C  11H  21O   4     G    300.00   4000.00 1384.00      1
 .426675367E+02 .481355870E-01-.164385340E-04 .254942818E-08-.147838407E-12    2
-.850035553E+05-.184014175E+03 .443641793E+01 .133210481E+00-.883606205E-04    3
 .302231077E-07-.426647212E-11-.712160785E+05 .229630078E+02                   4
QMDOOH                  C  11H  21O   4     G    300.00   4000.00 1378.00      1
 .463512360E+02 .442905004E-01-.156791241E-04 .249437540E-08-.147109263E-12    2
-.802179278E+05-.202701285E+03 .505901193E+01 .130586874E+00-.811966955E-04    3
 .236808295E-07-.254638441E-11-.648189073E+05 .227472201E+02                   4
ZMDOOH                  C  11H  21O   6     G    300.00   4000.00 1384.00      1
 .493171232E+02 .461887725E-01-.155948619E-04 .242596048E-08-.141314237E-12    2
-.997314376E+05-.213131636E+03 .613115269E+01 .145831804E+00-.103807590E-03    3
 .382530920E-07-.579145154E-11-.845666547E+05 .193222210E+02                   4
C12H7                   C  12H   7          G    300.00   4000.00 1000.00      1
 .119534365E+02 .523860720E-01-.276952580E-04 .698583900E-08-.684938540E-12    2
 .531995141E+05-.403925438E+02-.733802700E+01 .111965800E+00-.932829430E-04    3
 .358663430E-07-.426602200E-11 .580597660E+05 .573507160E+02                   4
RBIPHENYL               C  12H   9          G    300.00   4000.00 1000.00      1
 .214890352E+02 .375797860E-01-.121080230E-04 .129882780E-08 .000000000E+00    2
 .415521488E+05-.916763235E+02-.783196500E+01 .114327200E+00-.776398370E-04    3
 .194042280E-07 .000000000E+00 .498170300E+05 .608493300E+02                   4
NC12H25                 C  12H  25          G    300.00   4000.00 1387.00      1
 .379559371E+02 .541231481E-01-.184408520E-04 .285618139E-08-.165452331E-12    2
-.312698454E+05-.166157365E+03-.117025753E+01 .136564242E+00-.813840519E-04    3
 .231564976E-07-.240764498E-11-.167979250E+05 .471339366E+02                   4
NC12H25-OO              C  12H  25O   2     G    300.00   4000.00 1392.00      1
 .410672882E+02 .571682582E-01-.196096581E-04 .304996352E-08-.177163659E-12    2
-.498119415E+05-.176403781E+03 .761653139E+00 .147870053E+00-.980093227E-04    3
 .342486611E-07-.502171364E-11-.353144020E+05 .415448990E+02                   4
NC12-QOOH               C  12H  25O   2     G    300.00   4000.00 1392.00      1
 .427882927E+02 .547351985E-01-.185693137E-04 .286771608E-08-.165782124E-12    2
-.451897912E+05-.183774591E+03 .457142729E+00 .149660990E+00-.984019129E-04    3
 .327982507E-07-.438634589E-11-.301386488E+05 .448987214E+02                   4
NC12-OOQOOH             C  12H  25O   4     G    300.00   4000.00 1393.00      1
 .478223133E+02 .563342752E-01-.193784199E-04 .302016363E-08-.175696376E-12    2
-.648031378E+05-.208209874E+03 .250560092E+01 .157994999E+00-.105503812E-03    3
 .358709948E-07-.494871123E-11-.486270464E+05 .366890378E+02                   4
C14H9                   C  14H   9          G    300.00   4000.00 1000.00      1
 .255171870E+02 .393727940E-01-.123155080E-04 .127852800E-08 .000000000E+00    2
 .431324738E+05-.115618425E+03-.909474100E+01 .131333800E+00-.924017290E-04    3
 .240156710E-07 .000000000E+00 .527750200E+05 .639753600E+02                   4
C16H9                   C  16H   9          G    300.00   4000.00 1000.00      1
 .161628784E+02 .696969850E-01-.371786410E-04 .946306230E-08-.935417110E-12    2
 .461067047E+05-.652717249E+02-.114972670E+02 .151166960E+00-.116351410E-03    3
 .317097570E-07 .218082760E-11 .532378630E+05 .757195740E+02                   4
NC16H33                 C  16H  33          G    300.00   4000.00 1387.00      1
 .510324990E+02 .711045684E-01-.240491592E-04 .370710805E-08-.214054039E-12    2
-.477151440E+05-.228063103E+03-.243005348E+01 .186692969E+00-.115724867E-03    3
 .350879669E-07-.405848895E-11-.282942913E+05 .622394761E+02                   4
IC16H33                 C  16H  33          G    300.00   4000.00 1398.00      1
 .560389730E+02 .668182464E-01-.225681513E-04 .347608102E-08-.200620637E-12    2
-.583645424E+05-.270643351E+03-.953227198E+01 .224283987E+00-.166371012E-03    3
 .627848165E-07-.951119300E-11-.362947496E+05 .795385858E+02                   4
NC16-QOOH               C  16H  33O   2     G    300.00   4000.00 1394.00      1
 .557196631E+02 .758805933E-01-.260092776E-04 .404350192E-08-.234807139E-12    2
-.852319237E+05-.250905152E+03-.858601178E+00 .204663464E+00-.138309577E-03    3
 .488963438E-07-.717831502E-11-.651200924E+05 .543621098E+02                   4
IC16-QOOH               C  16H  33O   2     G    300.00   4000.00 1399.00      1
 .615798034E+02 .683372119E-01-.235040286E-04 .366308625E-08-.213104512E-12    2
-.710887760E+05-.294961987E+03-.836284759E+01 .243137667E+00-.193204766E-03    3
 .794478202E-07-.132585716E-10-.480052296E+05 .765156723E+02                   4
NC16H33-OO              C  16H  33O   2     G    300.00   4000.00 1392.00      1
 .537254976E+02 .751675700E-01-.257930312E-04 .401271756E-08-.233130903E-12    2
-.661992854E+05-.238675214E+03 .121036107E+00 .195526928E+00-.129332034E-03    3
 .448994551E-07-.651714304E-11-.469097176E+05 .512502917E+02                   4
IC16T-QOOH              C  16H  33O   2     G    300.00   4000.00 1397.00      1
 .619590914E+02 .670805941E-01-.228781110E-04 .354645272E-08-.205581639E-12    2
-.737750910E+05-.297686975E+03-.828638110E+01 .240615134E+00-.188046280E-03    3
 .753924180E-07-.122092604E-10-.505105835E+05 .759168895E+02                   4
IC16H33-OO              C  16H  33O   2     G    300.00   4000.00 1397.00      1
 .600009189E+02 .697612153E-01-.240119992E-04 .374399505E-08-.217877031E-12    2
-.771125672E+05-.288496873E+03-.807177622E+01 .238256241E+00-.186291159E-03    3
 .758296536E-07-.125956694E-10-.544214916E+05 .737310481E+02                   4
NC16-OOQOOH             C  16H  33O   4     G    300.00   4000.00 1393.00      1
 .605564321E+02 .743085731E-01-.255622121E-04 .398394439E-08-.231762903E-12    2
-.812450313E+05-.270973587E+03 .185761468E+01 .205470409E+00-.136236709E-03    3
 .460471713E-07-.632675050E-11-.602164277E+05 .464682670E+02                   4
IC16-OOQOOH             C  16H  33O   4     G    300.00   4000.00 1395.00      1
 .657312368E+02 .698159219E-01-.241818212E-04 .378635278E-08-.220988765E-12    2
-.891725518E+05-.313140345E+03-.709314164E+01 .252307521E+00-.202956898E-03    3
 .848048060E-07-.144255682E-10-.650715559E+05 .736645741E+02                   4
IC16T-OOQOOH            C  16H  33O   4     G    300.00   4000.00 1396.00      1
 .664600695E+02 .692200495E-01-.239811044E-04 .375550159E-08-.219211037E-12    2
-.927495777E+05-.318609160E+03-.734744585E+01 .256652224E+00-.210530384E-03    3
 .896944245E-07-.155165690E-10-.685533247E+05 .725686554E+02                   4
RUME16                  C  17H  31O   2     G    300.00   4000.00 1836.00      1
 .492312959E+02 .809629787E-01-.290414743E-04 .466984560E-08-.277987170E-12    2
-.712766099E+05-.212350222E+03 .581847898E+00 .197335153E+00-.132222747E-03    3
 .454132116E-07-.638160297E-11-.555076491E+05 .468001664E+02                   4
RMPAX                   C  17H  33O   2     G    300.00   4000.00 1000.00      1
 .347969412E+02 .108174887E+00-.436560662E-04 .805036686E-08-.557001848E-12    2
-.833532968E+05-.136711346E+03 .118429649E+02 .108281798E+00 .937470576E-04    3
-.175260710E-06 .681980157E-10-.741770519E+05-.304443036E+01                   4
QMPAOOH                 C  17H  33O   4     G    300.00   4000.00 1378.00      1
 .463512360E+02 .442905004E-01-.156791241E-04 .249437540E-08-.147109263E-12    2
-.802179278E+05-.202701285E+03 .505901193E+01 .130586874E+00-.811966955E-04    3
 .236808295E-07-.254638441E-11-.648189073E+05 .227472201E+02                   4
RMPAOOX                 C  17H  33O   4     G    300.00   4000.00 1384.00      1
 .426675367E+02 .481355870E-01-.164385340E-04 .254942818E-08-.147838407E-12    2
-.850035553E+05-.184014175E+03 .443641793E+01 .133210481E+00-.883606205E-04    3
 .302231077E-07-.426647212E-11-.712160785E+05 .229630078E+02                   4
ZMPAOOH                 C  17H  33O   6     G    300.00   4000.00 1384.00      1
 .493171232E+02 .461887725E-01-.155948619E-04 .242596048E-08-.141314237E-12    2
-.997314376E+05-.213131636E+03 .613115269E+01 .145831804E+00-.103807590E-03    3
 .382530920E-07-.579145154E-11-.845666547E+05 .193222210E+02                   4
RMLIN1X                 C  19H  31O   2     G    300.00   4000.00 1830.00      1
 .515951901E+02 .848982968E-01-.306132424E-04 .493978264E-08-.294767670E-12    2
-.437090861E+05-.222319284E+03-.124182769E+01 .210470141E+00-.141012967E-03    3
 .480938977E-07-.668889816E-11-.265018940E+05 .594297783E+02                   4
RMLIN1A                 C  19H  31O   2     G    300.00   4000.00 1830.00      1
 .515951901E+02 .848982968E-01-.306132424E-04 .493978264E-08-.294767670E-12    2
-.437090861E+05-.222319284E+03-.124182769E+01 .210470141E+00-.141012967E-03    3
 .480938977E-07-.668889816E-11-.265018940E+05 .594297783E+02                   4
RMLIN1OOX               C  19H  31O   4     G    300.00   4000.00 1854.00      1
 .566771062E+02 .848718923E-01-.306165992E-04 .494186779E-08-.294961213E-12    2
-.712260452E+05-.243221478E+03-.182318626E+01 .229267759E+00-.163619600E-03    3
 .597071790E-07-.884702825E-11-.526983896E+05 .668009912E+02                   4
QMLIN1OOX               C  19H  31O   4     G    300.00   4000.00 1859.00      1
 .597198037E+02 .825172318E-01-.298594827E-04 .482987333E-08-.288709215E-12    2
-.679692648E+05-.260058551E+03-.300959205E+01 .239625356E+00-.176824958E-03    3
 .662378545E-07-.999748235E-11-.483423909E+05 .715224170E+02                   4
ZMLIN1OOX               C  19H  31O   6     G    300.00   4000.00 1844.00      1
 .633953698E+02 .840133680E-01-.304696355E-04 .493592631E-08-.295352525E-12    2
-.861431583E+05-.275575442E+03 .377427203E+00 .239045319E+00-.172299424E-03    3
 .627369839E-07-.920510825E-11-.661691485E+05 .585014961E+02                   4
RMLINX                  C  19H  33O   2     G    300.00   4000.00 1386.00      1
 .611078575E+02 .762751735E-01-.262266430E-04 .408707626E-08-.237771674E-12    2
-.683962704E+05-.275956500E+03-.144781566E+01 .215019809E+00-.142192171E-03    3
 .476963895E-07-.649336150E-11-.458716461E+05 .627347784E+02                   4
RMLINA                  C  19H  33O   2     G    300.00   4000.00 1386.00      1
 .611078575E+02 .762751735E-01-.262266430E-04 .408707626E-08-.237771674E-12    2
-.683962704E+05-.275956500E+03-.144781566E+01 .215019809E+00-.142192171E-03    3
 .476963895E-07-.649336150E-11-.458716461E+05 .627347784E+02                   4
RMLINOOX                C  19H  33O   4     G    300.00   4000.00 1840.00      1
 .561396497E+02 .898573320E-01-.323076347E-04 .520295879E-08-.310043109E-12    2
-.835647272E+05-.240835194E+03 .146002415E+01 .221120424E+00-.149309126E-03    3
 .517229930E-07-.733489301E-11-.658774535E+05 .502873652E+02                   4
QMLINOOX                C  19H  33O   4     G    300.00   4000.00 1830.00      1
 .592334771E+02 .871071695E-01-.313329462E-04 .504827960E-08-.300945381E-12    2
-.780101129E+05-.256778117E+03-.383425349E+00 .231626065E+00-.160960610E-03    3
 .566395921E-07-.805109149E-11-.589322117E+05 .599912602E+02                   4
ZMLINOOX                C  19H  33O   6     G    300.00   4000.00 1183.00      1
 .601829822E+02 .877246704E-01-.308673874E-04 .490011538E-08-.289106438E-12    2
-.959756017E+05-.274111539E+03 .888177201E+00 .245491279E+00-.188867182E-03    3
 .756398491E-07-.122061299E-10-.781464330E+05 .361650421E+02                   4
RMEOLES                 C  19H  35O   2     G    300.00   4000.00 1386.00      1
 .617968812E+02 .797287018E-01-.272798012E-04 .423721781E-08-.245941529E-12    2
-.826622063E+05-.278715034E+03-.296860913E-01 .215538273E+00-.139084893E-03    3
 .453526106E-07-.596335185E-11-.602711250E+05 .564905254E+02                   4
RMEOLEA                 C  19H  35O   2     G    300.00   4000.00 1386.00      1
 .617968812E+02 .797287018E-01-.272798012E-04 .423721781E-08-.245941529E-12    2
-.826622063E+05-.278715034E+03-.296860913E-01 .215538273E+00-.139084893E-03    3
 .453526106E-07-.596335185E-11-.602711250E+05 .564905254E+02                   4
RMEOLEOOX               C  19H  35O   4     G    300.00   4000.00 1799.00      1
 .565118676E+02 .949710722E-01-.342666750E-04 .553134168E-08-.330143553E-12    2
-.121723087E+06-.240377715E+03 .312228984E+01 .215930145E+00-.133878272E-03    3
 .413627115E-07-.514696341E-11-.103763030E+06 .464356398E+02                   4
QMEOLEOOH               C  19H  35O   4     G    300.00   4000.00 1825.00      1
 .578903822E+02 .960618008E-01-.345783142E-04 .557312937E-08-.332293982E-12    2
-.145787244E+06-.248797880E+03-.121085721E+01 .236084007E+00-.157011163E-03    3
 .530523572E-07-.729693062E-11-.126516243E+06 .664772594E+02                   4
ZMEOLEOOX               C  19H  35O   6     G    300.00   4000.00 1175.00      1
 .558298346E+02 .101939581E+00-.350749088E-04 .548251413E-08-.319925836E-12    2
-.108843753E+06-.228788516E+03 .196924109E+01 .244903891E+00-.177892306E-03    3
 .692918136E-07-.110530115E-10-.926192007E+05 .531689573E+02                   4
RSTEAX                  C  19H  37O   2     G    300.00   4000.00 1000.00      1
 .410838828E+02 .116388491E+00-.460844475E-04 .839784976E-08-.576703150E-12    2
-.912925804E+05-.167019971E+03 .115570681E+02 .131479341E+00 .799583356E-04    3
-.171755777E-06 .679701047E-10-.799964069E+05 .174630364E+01                   4
RMSTEAOOX               C  19H  37O   4     G    300.00   4000.00 1384.00      1
 .294145201E+02 .809900030E-01-.261520592E-04 .393935978E-08-.226643615E-12    2
-.317656348E+05-.119394359E+03 .329283081E+01 .226000653E+00-.143515509E-03    3
 .442428385E-07-.517811632E-11-.232845416E+05 .214592368E+02                   4
QMSTEAOOH               C  19H  37O   4     G    300.00   4000.00 1378.00      1
 .297828900E+02 .771449164E-01-.253926493E-04 .388430700E-08-.225914471E-12    2
-.317651562E+05-.119207488E+03 .391542481E+01 .223377046E+00-.136351584E-03    3
 .377005603E-07-.345802861E-11-.232839019E+05 .214376580E+02                   4
ZMSTEAOOH               C  19H  37O   6     G    300.00   4000.00 1384.00      1
 .300794787E+02 .502955745E-01-.168090526E-04 .259970193E-08-.151164888E-12    2
-.397961494E+04-.130229963E+02 .598820430E+01 .157430576E+00-.110701951E-03    3
 .400055584E-07-.590540707E-11-.291813417E+04 .432758910E+01                   4
